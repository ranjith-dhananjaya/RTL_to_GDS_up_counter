VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO up_counter
  CLASS BLOCK ;
  FOREIGN up_counter ;
  ORIGIN 1.900 0.000 ;
  SIZE 115.800 BY 102.000 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 61.000 90.800 61.800 91.000 ;
        RECT 34.800 90.200 61.800 90.800 ;
        RECT 1.200 81.600 2.000 86.200 ;
        RECT 4.400 81.600 5.200 89.800 ;
        RECT 10.800 81.600 11.600 90.200 ;
        RECT 12.400 81.600 13.200 90.200 ;
        RECT 34.800 89.600 35.600 90.200 ;
        RECT 38.000 90.000 39.000 90.200 ;
        RECT 17.200 81.600 18.000 86.200 ;
        RECT 20.400 81.600 21.200 86.200 ;
        RECT 23.600 81.600 24.400 89.000 ;
        RECT 31.600 81.600 32.400 86.200 ;
        RECT 34.800 81.600 35.600 86.200 ;
        RECT 38.000 81.600 38.800 86.200 ;
        RECT 44.400 81.600 45.200 86.200 ;
        RECT 47.600 81.600 48.400 86.200 ;
        RECT 55.600 81.600 56.400 86.200 ;
        RECT 58.800 81.600 59.600 86.200 ;
        RECT 62.000 81.600 62.800 86.200 ;
        RECT 65.200 81.600 66.000 86.200 ;
        RECT 68.400 81.600 69.400 88.800 ;
        RECT 74.600 82.200 75.600 88.800 ;
        RECT 74.600 81.600 75.400 82.200 ;
        RECT 86.000 81.600 86.800 89.000 ;
        RECT 89.200 81.600 90.000 86.200 ;
        RECT 92.400 81.600 93.200 85.800 ;
        RECT 97.200 81.600 98.000 89.800 ;
        RECT 100.400 81.600 101.200 86.200 ;
        RECT 102.000 81.600 102.800 86.200 ;
        RECT 105.200 81.600 106.000 86.200 ;
        RECT 108.400 81.600 109.200 89.000 ;
        RECT 0.400 80.400 111.600 81.600 ;
        RECT 1.200 75.800 2.000 80.400 ;
        RECT 4.400 75.800 5.200 80.400 ;
        RECT 7.600 75.800 8.400 80.400 ;
        RECT 10.800 75.800 11.600 80.400 ;
        RECT 18.800 75.800 19.600 80.400 ;
        RECT 22.000 75.800 22.800 80.400 ;
        RECT 28.400 75.800 29.200 80.400 ;
        RECT 31.600 75.800 32.400 80.400 ;
        RECT 34.800 75.800 35.600 80.400 ;
        RECT 41.200 75.800 42.000 80.400 ;
        RECT 44.400 75.800 45.200 80.400 ;
        RECT 47.600 75.800 48.400 80.400 ;
        RECT 54.000 75.800 54.800 80.400 ;
        RECT 57.200 75.800 58.000 80.400 ;
        RECT 65.200 75.800 66.000 80.400 ;
        RECT 68.400 75.800 69.200 80.400 ;
        RECT 71.600 75.800 72.400 80.400 ;
        RECT 74.800 75.800 75.600 80.400 ;
        RECT 28.200 71.800 29.000 72.000 ;
        RECT 31.600 71.800 32.400 72.400 ;
        RECT 5.400 71.200 32.400 71.800 ;
        RECT 44.400 71.800 45.200 72.400 ;
        RECT 47.800 71.800 48.600 72.000 ;
        RECT 81.200 71.800 82.000 80.400 ;
        RECT 86.000 71.800 86.800 80.400 ;
        RECT 92.400 73.800 93.200 80.400 ;
        RECT 105.200 73.000 106.000 80.400 ;
        RECT 44.400 71.200 71.400 71.800 ;
        RECT 5.400 71.000 6.200 71.200 ;
        RECT 70.600 71.000 71.400 71.200 ;
        RECT 30.600 50.800 31.400 51.000 ;
        RECT 4.400 50.200 31.400 50.800 ;
        RECT 4.400 49.600 5.200 50.200 ;
        RECT 7.600 50.000 8.600 50.200 ;
        RECT 1.200 41.600 2.000 46.200 ;
        RECT 4.400 41.600 5.200 46.200 ;
        RECT 7.600 41.600 8.400 46.200 ;
        RECT 14.000 41.600 14.800 46.200 ;
        RECT 17.200 41.600 18.000 46.200 ;
        RECT 25.200 41.600 26.000 46.200 ;
        RECT 28.400 41.600 29.200 46.200 ;
        RECT 31.600 41.600 32.400 46.200 ;
        RECT 34.800 41.600 35.600 46.200 ;
        RECT 42.800 41.600 43.800 48.800 ;
        RECT 49.000 42.200 50.000 48.800 ;
        RECT 49.000 41.600 49.800 42.200 ;
        RECT 55.600 41.600 56.400 49.000 ;
        RECT 62.000 41.600 62.800 50.200 ;
        RECT 63.600 41.600 64.400 46.200 ;
        RECT 66.800 41.600 67.600 46.200 ;
        RECT 68.400 41.600 69.200 50.200 ;
        RECT 73.200 41.600 74.000 46.200 ;
        RECT 84.400 41.600 85.200 50.200 ;
        RECT 87.600 41.600 88.400 45.800 ;
        RECT 90.800 41.600 91.600 46.200 ;
        RECT 94.000 41.600 94.800 49.000 ;
        RECT 98.800 41.600 99.600 49.000 ;
        RECT 103.600 41.600 104.400 49.000 ;
        RECT 0.400 40.400 111.600 41.600 ;
        RECT 1.200 31.800 2.000 40.400 ;
        RECT 4.400 31.800 5.200 40.400 ;
        RECT 6.000 35.800 6.800 40.400 ;
        RECT 9.200 35.800 10.000 40.400 ;
        RECT 12.400 35.800 13.200 40.400 ;
        RECT 18.800 35.800 19.600 40.400 ;
        RECT 22.000 35.800 22.800 40.400 ;
        RECT 30.000 35.800 30.800 40.400 ;
        RECT 33.200 35.800 34.000 40.400 ;
        RECT 36.400 35.800 37.200 40.400 ;
        RECT 39.600 35.800 40.400 40.400 ;
        RECT 9.200 31.800 10.000 32.400 ;
        RECT 12.600 31.800 13.400 32.000 ;
        RECT 49.200 31.800 50.000 40.400 ;
        RECT 50.800 35.800 51.600 40.400 ;
        RECT 54.000 35.800 54.800 40.400 ;
        RECT 57.200 35.800 58.000 40.400 ;
        RECT 63.600 35.800 64.400 40.400 ;
        RECT 66.800 35.800 67.600 40.400 ;
        RECT 74.800 35.800 75.600 40.400 ;
        RECT 78.000 35.800 78.800 40.400 ;
        RECT 81.200 35.800 82.000 40.400 ;
        RECT 84.400 35.800 85.200 40.400 ;
        RECT 92.400 36.200 93.200 40.400 ;
        RECT 95.600 35.800 96.400 40.400 ;
        RECT 98.800 35.800 99.600 40.400 ;
        RECT 102.000 33.000 102.800 40.400 ;
        RECT 106.800 33.000 107.600 40.400 ;
        RECT 54.000 31.800 54.800 32.400 ;
        RECT 57.200 31.800 58.200 32.000 ;
        RECT 9.200 31.200 36.200 31.800 ;
        RECT 54.000 31.200 81.000 31.800 ;
        RECT 35.400 31.000 36.200 31.200 ;
        RECT 80.200 31.000 81.000 31.200 ;
        RECT 30.600 10.800 31.400 11.000 ;
        RECT 81.800 10.800 82.600 11.000 ;
        RECT 4.400 10.200 31.400 10.800 ;
        RECT 55.600 10.200 82.600 10.800 ;
        RECT 4.400 9.600 5.200 10.200 ;
        RECT 7.800 10.000 8.600 10.200 ;
        RECT 55.600 9.600 56.400 10.200 ;
        RECT 59.000 10.000 59.800 10.200 ;
        RECT 1.200 1.600 2.000 6.200 ;
        RECT 4.400 1.600 5.200 6.200 ;
        RECT 7.600 1.600 8.400 6.200 ;
        RECT 14.000 1.600 14.800 6.200 ;
        RECT 17.200 1.600 18.000 6.200 ;
        RECT 25.200 1.600 26.000 6.200 ;
        RECT 28.400 1.600 29.200 6.200 ;
        RECT 31.600 1.600 32.400 6.200 ;
        RECT 34.800 1.600 35.600 6.200 ;
        RECT 42.800 1.600 43.800 8.800 ;
        RECT 49.000 2.200 50.000 8.800 ;
        RECT 49.000 1.600 49.800 2.200 ;
        RECT 52.400 1.600 53.200 6.200 ;
        RECT 55.600 1.600 56.400 6.200 ;
        RECT 58.800 1.600 59.600 6.200 ;
        RECT 65.200 1.600 66.000 6.200 ;
        RECT 68.400 1.600 69.200 6.200 ;
        RECT 76.400 1.600 77.200 6.200 ;
        RECT 79.600 1.600 80.400 6.200 ;
        RECT 82.800 1.600 83.600 6.200 ;
        RECT 86.000 1.600 86.800 6.200 ;
        RECT 92.400 1.600 93.200 6.200 ;
        RECT 95.600 1.600 96.400 6.200 ;
        RECT 98.800 1.600 99.600 6.200 ;
        RECT 100.400 1.600 101.200 6.200 ;
        RECT 103.600 1.600 104.400 10.200 ;
        RECT 107.800 1.600 108.600 6.200 ;
        RECT 0.400 0.400 111.600 1.600 ;
      LAYER via1 ;
        RECT 38.000 85.400 38.800 86.200 ;
        RECT 35.000 80.600 35.800 81.400 ;
        RECT 36.400 80.600 37.200 81.400 ;
        RECT 37.800 80.600 38.600 81.400 ;
        RECT 31.600 77.600 32.400 78.400 ;
        RECT 44.400 77.600 45.200 78.400 ;
        RECT 31.600 71.600 32.400 72.400 ;
        RECT 44.400 71.600 45.200 72.400 ;
        RECT 7.600 43.600 8.400 44.400 ;
        RECT 35.000 40.600 35.800 41.400 ;
        RECT 36.400 40.600 37.200 41.400 ;
        RECT 37.800 40.600 38.600 41.400 ;
        RECT 9.200 37.600 10.000 38.400 ;
        RECT 9.200 31.600 10.000 32.400 ;
        RECT 57.200 31.200 58.000 32.000 ;
        RECT 4.400 3.600 5.200 4.400 ;
        RECT 55.600 3.600 56.400 4.400 ;
        RECT 35.000 0.600 35.800 1.400 ;
        RECT 36.400 0.600 37.200 1.400 ;
        RECT 37.800 0.600 38.600 1.400 ;
      LAYER metal2 ;
        RECT 38.000 90.000 38.800 90.800 ;
        RECT 38.100 86.200 38.700 90.000 ;
        RECT 38.000 85.400 38.800 86.200 ;
        RECT 34.400 80.600 39.200 81.400 ;
        RECT 31.600 77.600 32.400 78.400 ;
        RECT 44.400 77.600 45.200 78.400 ;
        RECT 31.700 72.400 32.300 77.600 ;
        RECT 44.500 72.400 45.100 77.600 ;
        RECT 31.600 71.600 32.400 72.400 ;
        RECT 44.400 71.600 45.200 72.400 ;
        RECT 7.600 50.000 8.400 50.800 ;
        RECT 7.700 44.400 8.300 50.000 ;
        RECT 7.600 43.600 8.400 44.400 ;
        RECT 34.400 40.600 39.200 41.400 ;
        RECT 9.200 37.600 10.000 38.400 ;
        RECT 9.300 32.400 9.900 37.600 ;
        RECT 57.200 35.800 58.000 36.600 ;
        RECT 9.200 31.600 10.000 32.400 ;
        RECT 57.300 32.000 57.900 35.800 ;
        RECT 57.200 31.200 58.000 32.000 ;
        RECT 4.400 9.600 5.200 10.400 ;
        RECT 55.600 9.600 56.400 10.400 ;
        RECT 4.500 4.400 5.100 9.600 ;
        RECT 55.700 4.400 56.300 9.600 ;
        RECT 4.400 3.600 5.200 4.400 ;
        RECT 55.600 3.600 56.400 4.400 ;
        RECT 34.400 0.600 39.200 1.400 ;
      LAYER via2 ;
        RECT 35.000 80.600 35.800 81.400 ;
        RECT 36.400 80.600 37.200 81.400 ;
        RECT 37.800 80.600 38.600 81.400 ;
        RECT 35.000 40.600 35.800 41.400 ;
        RECT 36.400 40.600 37.200 41.400 ;
        RECT 37.800 40.600 38.600 41.400 ;
        RECT 35.000 0.600 35.800 1.400 ;
        RECT 36.400 0.600 37.200 1.400 ;
        RECT 37.800 0.600 38.600 1.400 ;
      LAYER metal3 ;
        RECT 34.400 80.400 39.200 81.600 ;
        RECT 34.400 40.400 39.200 41.600 ;
        RECT 34.400 0.400 39.200 1.600 ;
      LAYER via3 ;
        RECT 34.800 80.600 35.600 81.400 ;
        RECT 36.400 80.600 37.200 81.400 ;
        RECT 38.000 80.600 38.800 81.400 ;
        RECT 34.800 40.600 35.600 41.400 ;
        RECT 36.400 40.600 37.200 41.400 ;
        RECT 38.000 40.600 38.800 41.400 ;
        RECT 34.800 0.600 35.600 1.400 ;
        RECT 36.400 0.600 37.200 1.400 ;
        RECT 38.000 0.600 38.800 1.400 ;
      LAYER metal4 ;
        RECT 34.400 0.000 39.200 102.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.400 100.400 111.600 101.600 ;
        RECT 3.800 96.000 4.600 100.400 ;
        RECT 7.600 97.800 8.400 100.400 ;
        RECT 10.800 97.800 11.600 100.400 ;
        RECT 12.400 97.800 13.200 100.400 ;
        RECT 15.600 97.800 16.400 100.400 ;
        RECT 17.200 95.800 18.000 100.400 ;
        RECT 23.600 95.800 24.400 100.400 ;
        RECT 34.800 95.800 35.600 100.400 ;
        RECT 44.400 97.800 45.200 100.400 ;
        RECT 47.600 97.800 48.400 100.400 ;
        RECT 58.800 95.800 59.600 100.400 ;
        RECT 65.200 97.800 66.000 100.400 ;
        RECT 68.400 96.400 69.400 100.400 ;
        RECT 74.600 99.800 75.400 100.400 ;
        RECT 74.600 96.400 75.600 99.800 ;
        RECT 82.800 97.800 83.600 100.400 ;
        RECT 87.000 95.800 87.800 100.400 ;
        RECT 89.200 93.800 90.000 100.400 ;
        RECT 97.800 96.000 98.600 100.400 ;
        RECT 105.200 95.800 106.000 100.400 ;
        RECT 108.400 95.800 109.200 100.400 ;
        RECT 1.200 61.600 2.000 64.200 ;
        RECT 7.600 61.600 8.400 66.200 ;
        RECT 18.800 61.600 19.600 64.200 ;
        RECT 22.000 61.600 22.800 64.200 ;
        RECT 31.600 61.600 32.400 66.200 ;
        RECT 44.400 61.600 45.200 66.200 ;
        RECT 54.000 61.600 54.800 64.200 ;
        RECT 57.200 61.600 58.000 64.200 ;
        RECT 68.400 61.600 69.200 66.200 ;
        RECT 74.800 61.600 75.600 64.200 ;
        RECT 81.200 61.600 82.000 64.200 ;
        RECT 84.400 61.600 85.200 64.200 ;
        RECT 86.000 61.600 86.800 64.200 ;
        RECT 89.200 61.600 90.000 64.200 ;
        RECT 92.400 61.600 93.200 64.200 ;
        RECT 95.600 61.600 96.400 63.800 ;
        RECT 105.200 61.600 106.000 66.200 ;
        RECT 0.400 60.400 111.600 61.600 ;
        RECT 4.400 55.800 5.200 60.400 ;
        RECT 14.000 57.800 14.800 60.400 ;
        RECT 17.200 57.800 18.000 60.400 ;
        RECT 28.400 55.800 29.200 60.400 ;
        RECT 34.800 57.800 35.600 60.400 ;
        RECT 42.800 56.400 43.800 60.400 ;
        RECT 49.000 59.800 49.800 60.400 ;
        RECT 49.000 56.400 50.000 59.800 ;
        RECT 52.400 57.800 53.200 60.400 ;
        RECT 56.600 55.800 57.400 60.400 ;
        RECT 58.800 57.800 59.600 60.400 ;
        RECT 62.000 57.800 62.800 60.400 ;
        RECT 66.800 55.800 67.600 60.400 ;
        RECT 68.400 57.800 69.200 60.400 ;
        RECT 71.600 57.800 72.400 60.400 ;
        RECT 73.200 57.800 74.000 60.400 ;
        RECT 81.200 57.800 82.000 60.400 ;
        RECT 84.400 57.800 85.200 60.400 ;
        RECT 90.800 53.800 91.600 60.400 ;
        RECT 94.000 55.800 94.800 60.400 ;
        RECT 98.800 55.800 99.600 60.400 ;
        RECT 103.600 55.800 104.400 60.400 ;
        RECT 1.200 21.600 2.000 26.200 ;
        RECT 4.400 21.600 5.200 26.200 ;
        RECT 9.200 21.600 10.000 26.200 ;
        RECT 18.800 21.600 19.600 24.200 ;
        RECT 22.000 21.600 22.800 24.200 ;
        RECT 33.200 21.600 34.000 26.200 ;
        RECT 39.600 21.600 40.400 24.200 ;
        RECT 46.000 21.600 46.800 24.200 ;
        RECT 49.200 21.600 50.000 24.200 ;
        RECT 54.000 21.600 54.800 26.200 ;
        RECT 63.600 21.600 64.400 24.200 ;
        RECT 66.800 21.600 67.600 24.200 ;
        RECT 78.000 21.600 78.800 26.200 ;
        RECT 84.400 21.600 85.200 24.200 ;
        RECT 95.600 21.600 96.400 28.200 ;
        RECT 98.800 21.600 99.600 24.200 ;
        RECT 102.000 21.600 102.800 26.200 ;
        RECT 106.800 21.600 107.600 26.200 ;
        RECT 0.400 20.400 111.600 21.600 ;
        RECT 4.400 15.800 5.200 20.400 ;
        RECT 14.000 17.800 14.800 20.400 ;
        RECT 17.200 17.800 18.000 20.400 ;
        RECT 28.400 15.800 29.200 20.400 ;
        RECT 34.800 17.800 35.600 20.400 ;
        RECT 42.800 16.400 43.800 20.400 ;
        RECT 49.000 19.800 49.800 20.400 ;
        RECT 49.000 16.400 50.000 19.800 ;
        RECT 55.600 15.800 56.400 20.400 ;
        RECT 65.200 17.800 66.000 20.400 ;
        RECT 68.400 17.800 69.200 20.400 ;
        RECT 79.600 15.800 80.400 20.400 ;
        RECT 86.000 17.800 86.800 20.400 ;
        RECT 92.400 17.800 93.200 20.400 ;
        RECT 98.800 15.800 99.600 20.400 ;
        RECT 100.400 17.800 101.200 20.400 ;
        RECT 105.200 16.600 106.000 20.400 ;
      LAYER via1 ;
        RECT 79.800 100.600 80.600 101.400 ;
        RECT 81.200 100.600 82.000 101.400 ;
        RECT 82.600 100.600 83.400 101.400 ;
        RECT 79.800 60.600 80.600 61.400 ;
        RECT 81.200 60.600 82.000 61.400 ;
        RECT 82.600 60.600 83.400 61.400 ;
        RECT 79.800 20.600 80.600 21.400 ;
        RECT 81.200 20.600 82.000 21.400 ;
        RECT 82.600 20.600 83.400 21.400 ;
      LAYER metal2 ;
        RECT 79.200 100.600 84.000 101.400 ;
        RECT 79.200 60.600 84.000 61.400 ;
        RECT 79.200 20.600 84.000 21.400 ;
      LAYER via2 ;
        RECT 79.800 100.600 80.600 101.400 ;
        RECT 81.200 100.600 82.000 101.400 ;
        RECT 82.600 100.600 83.400 101.400 ;
        RECT 79.800 60.600 80.600 61.400 ;
        RECT 81.200 60.600 82.000 61.400 ;
        RECT 82.600 60.600 83.400 61.400 ;
        RECT 79.800 20.600 80.600 21.400 ;
        RECT 81.200 20.600 82.000 21.400 ;
        RECT 82.600 20.600 83.400 21.400 ;
      LAYER metal3 ;
        RECT 79.200 100.400 84.000 101.600 ;
        RECT 79.200 60.400 84.000 61.600 ;
        RECT 79.200 20.400 84.000 21.600 ;
      LAYER via3 ;
        RECT 79.600 100.600 80.400 101.400 ;
        RECT 81.200 100.600 82.000 101.400 ;
        RECT 82.800 100.600 83.600 101.400 ;
        RECT 79.600 60.600 80.400 61.400 ;
        RECT 81.200 60.600 82.000 61.400 ;
        RECT 82.800 60.600 83.600 61.400 ;
        RECT 79.600 20.600 80.400 21.400 ;
        RECT 81.200 20.600 82.000 21.400 ;
        RECT 82.800 20.600 83.600 21.400 ;
      LAYER metal4 ;
        RECT 79.200 0.000 84.000 102.000 ;
    END
  END gnd
  PIN enable
    PORT
      LAYER metal1 ;
        RECT 10.800 95.600 11.600 97.200 ;
        RECT 1.200 91.600 2.000 94.400 ;
        RECT 17.200 93.600 18.000 95.200 ;
      LAYER metal2 ;
        RECT 10.800 95.600 11.600 96.400 ;
        RECT 1.200 91.600 2.000 92.400 ;
        RECT 1.300 90.400 1.900 91.600 ;
        RECT 10.900 90.400 11.500 95.600 ;
        RECT 17.200 93.600 18.000 94.400 ;
        RECT 17.300 90.400 17.900 93.600 ;
        RECT 1.200 89.600 2.000 90.400 ;
        RECT 10.800 89.600 11.600 90.400 ;
        RECT 17.200 89.600 18.000 90.400 ;
      LAYER metal3 ;
        RECT 1.200 90.300 2.000 90.400 ;
        RECT 10.800 90.300 11.600 90.400 ;
        RECT 17.200 90.300 18.000 90.400 ;
        RECT -1.900 89.700 18.000 90.300 ;
        RECT 1.200 89.600 2.000 89.700 ;
        RECT 10.800 89.600 11.600 89.700 ;
        RECT 17.200 89.600 18.000 89.700 ;
    END
  END enable
  PIN clk
    PORT
      LAYER metal1 ;
        RECT 47.600 95.600 49.200 96.400 ;
        RECT 18.000 65.600 19.600 66.400 ;
        RECT 57.200 65.600 58.800 66.400 ;
        RECT 17.200 55.600 18.800 56.400 ;
        RECT 22.000 25.600 23.600 26.400 ;
        RECT 66.800 25.600 68.400 26.400 ;
        RECT 17.200 15.600 18.800 16.400 ;
        RECT 68.400 15.600 70.000 16.400 ;
      LAYER via1 ;
        RECT 18.800 65.600 19.600 66.400 ;
      LAYER metal2 ;
        RECT 47.600 95.600 48.400 96.400 ;
        RECT 47.700 66.400 48.300 95.600 ;
        RECT 18.800 65.600 19.600 66.400 ;
        RECT 47.600 65.600 48.400 66.400 ;
        RECT 57.200 65.600 58.000 66.400 ;
        RECT 18.900 60.300 19.500 65.600 ;
        RECT 17.300 59.700 19.500 60.300 ;
        RECT 17.300 56.400 17.900 59.700 ;
        RECT 17.200 55.600 18.000 56.400 ;
        RECT 17.300 38.400 17.900 55.600 ;
        RECT 17.200 37.600 18.000 38.400 ;
        RECT 22.000 37.600 22.800 38.400 ;
        RECT 22.100 32.400 22.700 37.600 ;
        RECT 22.000 31.600 22.800 32.400 ;
        RECT 22.100 26.400 22.700 31.600 ;
        RECT 22.000 25.600 22.800 26.400 ;
        RECT 66.800 25.600 67.600 26.400 ;
        RECT 22.100 20.400 22.700 25.600 ;
        RECT 66.900 20.400 67.500 25.600 ;
        RECT 17.200 19.600 18.000 20.400 ;
        RECT 22.000 19.600 22.800 20.400 ;
        RECT 66.800 19.600 67.600 20.400 ;
        RECT 68.400 19.600 69.200 20.400 ;
        RECT 17.300 16.400 17.900 19.600 ;
        RECT 68.500 16.400 69.100 19.600 ;
        RECT 17.200 15.600 18.000 16.400 ;
        RECT 68.400 15.600 69.200 16.400 ;
      LAYER metal3 ;
        RECT 18.800 66.300 19.600 66.400 ;
        RECT 47.600 66.300 48.400 66.400 ;
        RECT 57.200 66.300 58.000 66.400 ;
        RECT 18.800 65.700 58.000 66.300 ;
        RECT 18.800 65.600 19.600 65.700 ;
        RECT 47.600 65.600 48.400 65.700 ;
        RECT 57.200 65.600 58.000 65.700 ;
        RECT 17.200 38.300 18.000 38.400 ;
        RECT 22.000 38.300 22.800 38.400 ;
        RECT 17.200 37.700 22.800 38.300 ;
        RECT 17.200 37.600 18.000 37.700 ;
        RECT 22.000 37.600 22.800 37.700 ;
        RECT 22.000 32.300 22.800 32.400 ;
        RECT -1.900 31.700 22.800 32.300 ;
        RECT 22.000 31.600 22.800 31.700 ;
        RECT 17.200 20.300 18.000 20.400 ;
        RECT 22.000 20.300 22.800 20.400 ;
        RECT 66.800 20.300 67.600 20.400 ;
        RECT 68.400 20.300 69.200 20.400 ;
        RECT 17.200 19.700 69.200 20.300 ;
        RECT 17.200 19.600 18.000 19.700 ;
        RECT 22.000 19.600 22.800 19.700 ;
        RECT 66.800 19.600 67.600 19.700 ;
        RECT 68.400 19.600 69.200 19.700 ;
    END
  END clk
  PIN reset
    PORT
      LAYER metal1 ;
        RECT 1.200 26.800 2.000 28.400 ;
      LAYER via1 ;
        RECT 1.200 27.600 2.000 28.400 ;
      LAYER metal2 ;
        RECT 1.200 27.600 2.000 28.400 ;
      LAYER metal3 ;
        RECT 1.200 28.300 2.000 28.400 ;
        RECT -1.900 27.700 2.000 28.300 ;
        RECT 1.200 27.600 2.000 27.700 ;
    END
  END reset
  PIN out0
    PORT
      LAYER metal1 ;
        RECT 25.200 98.300 26.000 99.800 ;
        RECT 30.000 98.300 30.800 98.400 ;
        RECT 25.200 97.700 30.800 98.300 ;
        RECT 25.200 92.400 26.000 97.700 ;
        RECT 30.000 97.600 30.800 97.700 ;
        RECT 25.400 90.200 26.000 92.400 ;
        RECT 25.200 82.200 26.000 90.200 ;
      LAYER metal2 ;
        RECT 30.000 97.600 30.800 98.400 ;
      LAYER metal3 ;
        RECT 30.000 98.300 30.800 98.400 ;
        RECT 30.000 97.700 113.900 98.300 ;
        RECT 30.000 97.600 30.800 97.700 ;
    END
  END out0
  PIN out1
    PORT
      LAYER metal1 ;
        RECT 105.200 58.300 106.000 59.800 ;
        RECT 108.400 58.300 109.200 58.400 ;
        RECT 105.200 57.700 109.200 58.300 ;
        RECT 105.200 52.400 106.000 57.700 ;
        RECT 108.400 57.600 109.200 57.700 ;
        RECT 105.400 50.200 106.000 52.400 ;
        RECT 105.200 42.200 106.000 50.200 ;
      LAYER metal2 ;
        RECT 108.400 93.600 109.200 94.400 ;
        RECT 108.500 58.400 109.100 93.600 ;
        RECT 108.400 57.600 109.200 58.400 ;
      LAYER metal3 ;
        RECT 108.400 94.300 109.200 94.400 ;
        RECT 108.400 93.700 113.900 94.300 ;
        RECT 108.400 93.600 109.200 93.700 ;
    END
  END out1
  PIN out2
    PORT
      LAYER metal1 ;
        RECT 110.000 92.400 110.800 99.800 ;
        RECT 110.200 90.200 110.800 92.400 ;
        RECT 110.000 82.200 110.800 90.200 ;
      LAYER via1 ;
        RECT 110.000 87.600 110.800 88.400 ;
      LAYER metal2 ;
        RECT 110.000 89.600 110.800 90.400 ;
        RECT 110.100 88.400 110.700 89.600 ;
        RECT 110.000 87.600 110.800 88.400 ;
      LAYER metal3 ;
        RECT 110.000 90.300 110.800 90.400 ;
        RECT 110.000 89.700 113.900 90.300 ;
        RECT 110.000 89.600 110.800 89.700 ;
    END
  END out2
  PIN out3
    PORT
      LAYER metal1 ;
        RECT 106.800 71.800 107.600 79.800 ;
        RECT 107.000 69.600 107.600 71.800 ;
        RECT 106.800 68.300 107.600 69.600 ;
        RECT 110.000 68.300 110.800 68.400 ;
        RECT 106.800 67.700 110.800 68.300 ;
        RECT 106.800 62.200 107.600 67.700 ;
        RECT 110.000 67.600 110.800 67.700 ;
      LAYER metal2 ;
        RECT 110.000 69.600 110.800 70.400 ;
        RECT 110.100 68.400 110.700 69.600 ;
        RECT 110.000 67.600 110.800 68.400 ;
      LAYER metal3 ;
        RECT 110.000 70.300 110.800 70.400 ;
        RECT 110.000 69.700 113.900 70.300 ;
        RECT 110.000 69.600 110.800 69.700 ;
    END
  END out3
  PIN out4
    PORT
      LAYER metal1 ;
        RECT 100.400 52.400 101.200 59.800 ;
        RECT 100.600 50.200 101.200 52.400 ;
        RECT 100.400 42.200 101.200 50.200 ;
      LAYER via1 ;
        RECT 100.400 53.600 101.200 54.400 ;
      LAYER metal2 ;
        RECT 100.400 53.600 101.200 54.400 ;
      LAYER metal3 ;
        RECT 100.400 54.300 101.200 54.400 ;
        RECT 100.400 53.700 113.900 54.300 ;
        RECT 100.400 53.600 101.200 53.700 ;
    END
  END out4
  PIN out5
    PORT
      LAYER metal1 ;
        RECT 95.600 52.400 96.400 59.800 ;
        RECT 95.800 50.200 96.400 52.400 ;
        RECT 95.600 42.200 96.400 50.200 ;
      LAYER via1 ;
        RECT 95.600 47.600 96.400 48.400 ;
      LAYER metal2 ;
        RECT 95.600 49.600 96.400 50.400 ;
        RECT 95.700 48.400 96.300 49.600 ;
        RECT 95.600 47.600 96.400 48.400 ;
      LAYER metal3 ;
        RECT 95.600 50.300 96.400 50.400 ;
        RECT 95.600 49.700 113.900 50.300 ;
        RECT 95.600 49.600 96.400 49.700 ;
    END
  END out5
  PIN out6
    PORT
      LAYER metal1 ;
        RECT 103.600 31.800 104.400 39.800 ;
        RECT 103.800 29.600 104.400 31.800 ;
        RECT 103.600 22.200 104.400 29.600 ;
      LAYER via1 ;
        RECT 103.600 33.600 104.400 34.400 ;
      LAYER metal2 ;
        RECT 103.600 33.600 104.400 34.400 ;
      LAYER metal3 ;
        RECT 103.600 34.300 104.400 34.400 ;
        RECT 103.600 33.700 113.900 34.300 ;
        RECT 103.600 33.600 104.400 33.700 ;
    END
  END out6
  PIN out7
    PORT
      LAYER metal1 ;
        RECT 108.400 31.800 109.200 39.800 ;
        RECT 108.600 29.600 109.200 31.800 ;
        RECT 108.400 28.300 109.200 29.600 ;
        RECT 110.000 28.300 110.800 28.400 ;
        RECT 108.400 27.700 110.800 28.300 ;
        RECT 108.400 22.200 109.200 27.700 ;
        RECT 110.000 27.600 110.800 27.700 ;
      LAYER metal2 ;
        RECT 110.000 29.600 110.800 30.400 ;
        RECT 110.100 28.400 110.700 29.600 ;
        RECT 110.000 27.600 110.800 28.400 ;
      LAYER metal3 ;
        RECT 110.000 30.300 110.800 30.400 ;
        RECT 110.000 29.700 113.900 30.300 ;
        RECT 110.000 29.600 110.800 29.700 ;
    END
  END out7
  OBS
      LAYER metal1 ;
        RECT 1.200 95.800 2.000 99.800 ;
        RECT 5.400 96.800 6.200 99.800 ;
        RECT 9.200 97.800 10.000 99.800 ;
        RECT 14.000 97.800 14.800 99.800 ;
        RECT 5.400 95.800 6.800 96.800 ;
        RECT 1.400 95.600 2.000 95.800 ;
        RECT 1.400 95.200 3.200 95.600 ;
        RECT 1.400 95.000 5.600 95.200 ;
        RECT 2.600 94.600 5.600 95.000 ;
        RECT 4.800 94.400 5.600 94.600 ;
        RECT 3.200 93.800 4.000 94.000 ;
        RECT 3.000 93.200 4.000 93.800 ;
        RECT 3.000 92.400 3.600 93.200 ;
        RECT 2.800 91.600 3.600 92.400 ;
        RECT 4.800 91.000 5.400 94.400 ;
        RECT 6.200 92.400 6.800 95.800 ;
        RECT 9.200 94.400 9.800 97.800 ;
        RECT 12.400 95.600 13.200 97.200 ;
        RECT 9.200 94.300 10.000 94.400 ;
        RECT 12.500 94.300 13.100 95.600 ;
        RECT 14.200 94.400 14.800 97.800 ;
        RECT 19.800 96.400 20.600 99.800 ;
        RECT 9.200 93.700 13.100 94.300 ;
        RECT 9.200 93.600 10.000 93.700 ;
        RECT 14.000 93.600 14.800 94.400 ;
        RECT 6.000 91.600 6.800 92.400 ;
        RECT 3.000 90.400 5.400 91.000 ;
        RECT 3.000 86.200 3.600 90.400 ;
        RECT 6.200 90.200 6.800 91.600 ;
        RECT 7.600 90.800 8.400 92.400 ;
        RECT 9.200 90.200 9.800 93.600 ;
        RECT 14.200 90.200 14.800 93.600 ;
        RECT 18.800 95.600 21.200 96.400 ;
        RECT 15.600 90.800 16.400 92.400 ;
        RECT 2.800 82.200 3.600 86.200 ;
        RECT 6.000 82.200 6.800 90.200 ;
        RECT 8.200 89.400 10.000 90.200 ;
        RECT 14.000 89.400 15.800 90.200 ;
        RECT 8.200 82.200 9.000 89.400 ;
        RECT 15.000 84.400 15.800 89.400 ;
        RECT 15.000 83.600 16.400 84.400 ;
        RECT 15.000 82.200 15.800 83.600 ;
        RECT 18.800 82.200 19.600 95.600 ;
        RECT 22.000 95.200 22.800 99.800 ;
        RECT 22.000 94.600 24.200 95.200 ;
        RECT 22.000 92.300 22.800 93.200 ;
        RECT 20.500 91.700 22.800 92.300 ;
        RECT 20.500 90.400 21.100 91.700 ;
        RECT 22.000 91.600 22.800 91.700 ;
        RECT 23.600 91.600 24.200 94.600 ;
        RECT 31.600 93.800 32.400 99.800 ;
        RECT 38.000 96.600 38.800 99.800 ;
        RECT 39.600 97.000 40.400 99.800 ;
        RECT 41.200 97.000 42.000 99.800 ;
        RECT 42.800 97.000 43.600 99.800 ;
        RECT 46.000 97.000 46.800 99.800 ;
        RECT 49.200 97.000 50.000 99.800 ;
        RECT 50.800 97.000 51.600 99.800 ;
        RECT 52.400 97.000 53.200 99.800 ;
        RECT 54.000 97.000 54.800 99.800 ;
        RECT 36.200 95.800 38.800 96.600 ;
        RECT 55.600 96.600 56.400 99.800 ;
        RECT 42.200 95.800 46.800 96.400 ;
        RECT 36.200 95.200 37.000 95.800 ;
        RECT 34.000 94.400 37.000 95.200 ;
        RECT 31.600 93.000 40.400 93.800 ;
        RECT 42.200 93.400 43.000 95.800 ;
        RECT 46.000 95.600 46.800 95.800 ;
        RECT 52.200 95.600 53.200 96.400 ;
        RECT 55.600 95.800 58.000 96.600 ;
        RECT 44.400 93.600 45.200 95.200 ;
        RECT 46.000 94.800 46.800 95.000 ;
        RECT 46.000 94.200 50.400 94.800 ;
        RECT 49.600 94.000 50.400 94.200 ;
        RECT 23.600 90.800 24.800 91.600 ;
        RECT 20.400 88.800 21.200 90.400 ;
        RECT 23.600 90.200 24.200 90.800 ;
        RECT 22.000 89.600 24.200 90.200 ;
        RECT 22.000 82.200 22.800 89.600 ;
        RECT 31.600 87.400 32.400 93.000 ;
        RECT 41.000 92.600 43.000 93.400 ;
        RECT 46.800 92.600 50.000 93.400 ;
        RECT 52.400 92.800 53.200 95.600 ;
        RECT 57.200 95.200 58.000 95.800 ;
        RECT 57.200 94.600 59.000 95.200 ;
        RECT 58.200 93.400 59.000 94.600 ;
        RECT 62.000 94.600 62.800 99.800 ;
        RECT 63.600 96.000 64.400 99.800 ;
        RECT 63.600 95.200 64.600 96.000 ;
        RECT 66.800 95.800 67.600 99.800 ;
        RECT 71.200 96.200 72.800 99.800 ;
        RECT 66.800 95.200 69.200 95.800 ;
        RECT 62.000 94.000 63.200 94.600 ;
        RECT 58.200 92.600 62.000 93.400 ;
        RECT 33.000 92.000 33.800 92.200 ;
        RECT 38.000 92.000 38.800 92.400 ;
        RECT 55.600 92.000 56.400 92.600 ;
        RECT 62.600 92.000 63.200 94.000 ;
        RECT 33.000 91.400 56.400 92.000 ;
        RECT 62.400 91.400 63.200 92.000 ;
        RECT 63.800 94.300 64.600 95.200 ;
        RECT 68.400 95.000 69.200 95.200 ;
        RECT 69.800 94.800 70.600 95.600 ;
        RECT 69.800 94.400 70.400 94.800 ;
        RECT 66.800 94.300 68.400 94.400 ;
        RECT 63.800 93.700 68.400 94.300 ;
        RECT 62.400 89.600 63.000 91.400 ;
        RECT 63.800 90.800 64.600 93.700 ;
        RECT 66.800 93.600 68.400 93.700 ;
        RECT 69.600 93.600 70.400 94.400 ;
        RECT 71.200 92.800 71.800 96.200 ;
        RECT 76.400 95.800 77.200 99.800 ;
        RECT 83.000 96.400 83.800 97.200 ;
        RECT 72.400 95.400 74.000 95.600 ;
        RECT 72.400 94.800 74.400 95.400 ;
        RECT 75.000 95.200 77.200 95.800 ;
        RECT 82.800 95.600 83.600 96.400 ;
        RECT 84.400 95.800 85.200 99.800 ;
        RECT 75.000 95.000 75.800 95.200 ;
        RECT 73.800 94.400 74.400 94.800 ;
        RECT 72.400 93.400 73.200 94.200 ;
        RECT 73.800 93.800 77.200 94.400 ;
        RECT 75.600 93.600 77.200 93.800 ;
        RECT 70.800 92.400 71.800 92.800 ;
        RECT 65.200 92.300 66.000 92.400 ;
        RECT 70.000 92.300 71.800 92.400 ;
        RECT 65.200 92.200 71.800 92.300 ;
        RECT 72.600 92.800 73.200 93.400 ;
        RECT 72.600 92.200 75.200 92.800 ;
        RECT 65.200 91.700 71.400 92.200 ;
        RECT 74.400 92.000 75.200 92.200 ;
        RECT 82.800 92.200 83.600 92.400 ;
        RECT 84.600 92.200 85.200 95.800 ;
        RECT 86.000 92.800 86.800 94.400 ;
        RECT 92.800 94.200 93.600 99.800 ;
        RECT 96.200 96.800 97.000 99.800 ;
        RECT 95.600 95.800 97.000 96.800 ;
        RECT 100.400 95.800 101.200 99.800 ;
        RECT 102.600 96.400 103.400 99.800 ;
        RECT 102.600 95.800 104.400 96.400 ;
        RECT 92.800 93.800 94.600 94.200 ;
        RECT 93.000 93.600 94.600 93.800 ;
        RECT 87.600 92.200 88.400 92.400 ;
        RECT 65.200 91.600 66.000 91.700 ;
        RECT 70.000 91.600 71.400 91.700 ;
        RECT 82.800 91.600 85.200 92.200 ;
        RECT 86.800 91.600 88.400 92.200 ;
        RECT 90.800 91.600 92.400 92.400 ;
        RECT 41.200 89.400 42.000 89.600 ;
        RECT 36.600 89.000 42.000 89.400 ;
        RECT 35.800 88.800 42.000 89.000 ;
        RECT 43.000 89.000 51.600 89.600 ;
        RECT 33.200 88.000 34.800 88.800 ;
        RECT 35.800 88.200 37.200 88.800 ;
        RECT 43.000 88.200 43.600 89.000 ;
        RECT 50.800 88.800 51.600 89.000 ;
        RECT 54.000 89.000 63.000 89.600 ;
        RECT 54.000 88.800 54.800 89.000 ;
        RECT 34.200 87.600 34.800 88.000 ;
        RECT 37.800 87.600 43.600 88.200 ;
        RECT 44.200 87.600 46.800 88.400 ;
        RECT 31.600 86.800 33.600 87.400 ;
        RECT 34.200 86.800 38.400 87.600 ;
        RECT 33.000 86.200 33.600 86.800 ;
        RECT 33.000 85.600 34.000 86.200 ;
        RECT 33.200 82.200 34.000 85.600 ;
        RECT 36.400 82.200 37.200 86.800 ;
        RECT 39.600 82.200 40.400 85.000 ;
        RECT 41.200 82.200 42.000 85.000 ;
        RECT 42.800 82.200 43.600 87.000 ;
        RECT 46.000 82.200 46.800 87.000 ;
        RECT 49.200 82.200 50.000 88.400 ;
        RECT 57.200 87.600 59.800 88.400 ;
        RECT 52.400 86.800 56.600 87.600 ;
        RECT 50.800 82.200 51.600 85.000 ;
        RECT 52.400 82.200 53.200 85.000 ;
        RECT 54.000 82.200 54.800 85.000 ;
        RECT 57.200 82.200 58.000 87.600 ;
        RECT 62.400 87.400 63.000 89.000 ;
        RECT 60.400 86.800 63.000 87.400 ;
        RECT 63.600 90.000 64.600 90.800 ;
        RECT 70.800 90.200 71.400 91.600 ;
        RECT 72.200 91.400 73.000 91.600 ;
        RECT 72.200 90.800 75.600 91.400 ;
        RECT 75.000 90.200 75.600 90.800 ;
        RECT 83.000 90.200 83.600 91.600 ;
        RECT 86.800 91.200 87.600 91.600 ;
        RECT 89.200 90.300 90.000 91.200 ;
        RECT 94.000 90.400 94.600 93.600 ;
        RECT 95.600 92.400 96.200 95.800 ;
        RECT 100.400 95.600 101.000 95.800 ;
        RECT 99.200 95.200 101.000 95.600 ;
        RECT 96.800 95.000 101.000 95.200 ;
        RECT 96.800 94.600 99.800 95.000 ;
        RECT 96.800 94.400 97.600 94.600 ;
        RECT 95.600 91.600 96.400 92.400 ;
        RECT 90.800 90.300 91.600 90.400 ;
        RECT 60.400 82.200 61.200 86.800 ;
        RECT 63.600 82.200 64.400 90.000 ;
        RECT 66.800 89.600 69.200 90.200 ;
        RECT 70.800 89.600 72.800 90.200 ;
        RECT 66.800 82.200 67.600 89.600 ;
        RECT 68.400 89.400 69.200 89.600 ;
        RECT 71.200 82.200 72.800 89.600 ;
        RECT 75.000 89.600 77.200 90.200 ;
        RECT 75.000 89.400 75.800 89.600 ;
        RECT 76.400 82.200 77.200 89.600 ;
        RECT 81.200 84.300 82.000 84.400 ;
        RECT 82.800 84.300 83.600 90.200 ;
        RECT 81.200 83.700 83.600 84.300 ;
        RECT 81.200 83.600 82.000 83.700 ;
        RECT 82.800 82.200 83.600 83.700 ;
        RECT 84.400 89.600 88.400 90.200 ;
        RECT 89.200 89.700 91.600 90.300 ;
        RECT 89.200 89.600 90.000 89.700 ;
        RECT 90.800 89.600 91.600 89.700 ;
        RECT 94.000 89.600 94.800 90.400 ;
        RECT 95.600 90.200 96.200 91.600 ;
        RECT 97.000 91.000 97.600 94.400 ;
        RECT 98.400 93.800 99.200 94.000 ;
        RECT 98.400 93.200 99.400 93.800 ;
        RECT 98.800 92.400 99.400 93.200 ;
        RECT 100.400 92.800 101.200 94.400 ;
        RECT 98.800 91.600 99.600 92.400 ;
        RECT 97.000 90.400 99.400 91.000 ;
        RECT 84.400 82.200 85.200 89.600 ;
        RECT 87.600 82.200 88.400 89.600 ;
        RECT 92.400 87.600 93.200 89.200 ;
        RECT 94.000 87.000 94.600 89.600 ;
        RECT 91.000 86.400 94.600 87.000 ;
        RECT 91.000 86.200 91.600 86.400 ;
        RECT 90.800 82.200 91.600 86.200 ;
        RECT 94.000 86.200 94.600 86.400 ;
        RECT 94.000 82.200 94.800 86.200 ;
        RECT 95.600 82.200 96.400 90.200 ;
        RECT 98.800 86.200 99.400 90.400 ;
        RECT 102.000 88.800 102.800 90.400 ;
        RECT 98.800 82.200 99.600 86.200 ;
        RECT 103.600 82.200 104.400 95.800 ;
        RECT 106.800 95.200 107.600 99.800 ;
        RECT 105.200 93.600 106.000 95.200 ;
        RECT 106.800 94.600 109.000 95.200 ;
        RECT 106.800 91.600 107.600 93.200 ;
        RECT 108.400 91.600 109.000 94.600 ;
        RECT 108.400 90.800 109.600 91.600 ;
        RECT 108.400 90.200 109.000 90.800 ;
        RECT 106.800 89.600 109.000 90.200 ;
        RECT 106.800 82.200 107.600 89.600 ;
        RECT 2.800 72.000 3.600 79.800 ;
        RECT 6.000 75.200 6.800 79.800 ;
        RECT 2.600 71.200 3.600 72.000 ;
        RECT 4.200 74.600 6.800 75.200 ;
        RECT 4.200 73.000 4.800 74.600 ;
        RECT 9.200 74.400 10.000 79.800 ;
        RECT 12.400 77.000 13.200 79.800 ;
        RECT 14.000 77.000 14.800 79.800 ;
        RECT 15.600 77.000 16.400 79.800 ;
        RECT 10.600 74.400 14.800 75.200 ;
        RECT 7.400 73.600 10.000 74.400 ;
        RECT 17.200 73.600 18.000 79.800 ;
        RECT 20.400 75.000 21.200 79.800 ;
        RECT 23.600 75.000 24.400 79.800 ;
        RECT 25.200 77.000 26.000 79.800 ;
        RECT 26.800 77.000 27.600 79.800 ;
        RECT 30.000 75.200 30.800 79.800 ;
        RECT 33.200 76.400 34.000 79.800 ;
        RECT 42.800 76.400 43.600 79.800 ;
        RECT 33.200 75.800 34.200 76.400 ;
        RECT 33.600 75.200 34.200 75.800 ;
        RECT 42.600 75.800 43.600 76.400 ;
        RECT 42.600 75.200 43.200 75.800 ;
        RECT 46.000 75.200 46.800 79.800 ;
        RECT 49.200 77.000 50.000 79.800 ;
        RECT 50.800 77.000 51.600 79.800 ;
        RECT 28.800 74.400 33.000 75.200 ;
        RECT 33.600 74.600 35.600 75.200 ;
        RECT 20.400 73.600 23.000 74.400 ;
        RECT 23.600 73.800 29.400 74.400 ;
        RECT 32.400 74.000 33.000 74.400 ;
        RECT 12.400 73.000 13.200 73.200 ;
        RECT 4.200 72.400 13.200 73.000 ;
        RECT 15.600 73.000 16.400 73.200 ;
        RECT 23.600 73.000 24.200 73.800 ;
        RECT 30.000 73.200 31.400 73.800 ;
        RECT 32.400 73.200 34.000 74.000 ;
        RECT 15.600 72.400 24.200 73.000 ;
        RECT 25.200 73.000 31.400 73.200 ;
        RECT 25.200 72.600 30.600 73.000 ;
        RECT 25.200 72.400 26.000 72.600 ;
        RECT 2.600 66.800 3.400 71.200 ;
        RECT 4.200 70.600 4.800 72.400 ;
        RECT 4.000 70.000 4.800 70.600 ;
        RECT 10.800 70.000 34.200 70.600 ;
        RECT 4.000 68.000 4.600 70.000 ;
        RECT 10.800 69.400 11.600 70.000 ;
        RECT 28.400 69.600 29.200 70.000 ;
        RECT 33.200 69.800 34.200 70.000 ;
        RECT 33.200 69.600 34.000 69.800 ;
        RECT 5.200 68.600 9.000 69.400 ;
        RECT 4.000 67.400 5.200 68.000 ;
        RECT 2.600 66.000 3.600 66.800 ;
        RECT 2.800 62.200 3.600 66.000 ;
        RECT 4.400 62.200 5.200 67.400 ;
        RECT 8.200 67.400 9.000 68.600 ;
        RECT 8.200 66.800 10.000 67.400 ;
        RECT 9.200 66.200 10.000 66.800 ;
        RECT 14.000 66.400 14.800 69.200 ;
        RECT 17.200 68.600 20.400 69.400 ;
        RECT 24.200 68.600 26.200 69.400 ;
        RECT 34.800 69.000 35.600 74.600 ;
        RECT 16.800 67.800 17.600 68.000 ;
        RECT 16.800 67.200 21.200 67.800 ;
        RECT 20.400 67.000 21.200 67.200 ;
        RECT 22.000 66.800 22.800 68.400 ;
        RECT 9.200 65.400 11.600 66.200 ;
        RECT 14.000 65.600 15.000 66.400 ;
        RECT 20.400 66.200 21.200 66.400 ;
        RECT 24.200 66.200 25.000 68.600 ;
        RECT 26.800 68.200 35.600 69.000 ;
        RECT 30.200 66.800 33.200 67.600 ;
        RECT 30.200 66.200 31.000 66.800 ;
        RECT 20.400 65.600 25.000 66.200 ;
        RECT 10.800 62.200 11.600 65.400 ;
        RECT 28.400 65.400 31.000 66.200 ;
        RECT 12.400 62.200 13.200 65.000 ;
        RECT 14.000 62.200 14.800 65.000 ;
        RECT 15.600 62.200 16.400 65.000 ;
        RECT 17.200 62.200 18.000 65.000 ;
        RECT 20.400 62.200 21.200 65.000 ;
        RECT 23.600 62.200 24.400 65.000 ;
        RECT 25.200 62.200 26.000 65.000 ;
        RECT 26.800 62.200 27.600 65.000 ;
        RECT 28.400 62.200 29.200 65.400 ;
        RECT 34.800 62.200 35.600 68.200 ;
        RECT 41.200 74.600 43.200 75.200 ;
        RECT 41.200 69.000 42.000 74.600 ;
        RECT 43.800 74.400 48.000 75.200 ;
        RECT 52.400 75.000 53.200 79.800 ;
        RECT 55.600 75.000 56.400 79.800 ;
        RECT 43.800 74.000 44.400 74.400 ;
        RECT 42.800 73.200 44.400 74.000 ;
        RECT 47.400 73.800 53.200 74.400 ;
        RECT 45.400 73.200 46.800 73.800 ;
        RECT 45.400 73.000 51.600 73.200 ;
        RECT 46.200 72.600 51.600 73.000 ;
        RECT 50.800 72.400 51.600 72.600 ;
        RECT 52.600 73.000 53.200 73.800 ;
        RECT 53.800 73.600 56.400 74.400 ;
        RECT 58.800 73.600 59.600 79.800 ;
        RECT 60.400 77.000 61.200 79.800 ;
        RECT 62.000 77.000 62.800 79.800 ;
        RECT 63.600 77.000 64.400 79.800 ;
        RECT 62.000 74.400 66.200 75.200 ;
        RECT 66.800 74.400 67.600 79.800 ;
        RECT 70.000 75.200 70.800 79.800 ;
        RECT 70.000 74.600 72.600 75.200 ;
        RECT 66.800 73.600 69.400 74.400 ;
        RECT 60.400 73.000 61.200 73.200 ;
        RECT 52.600 72.400 61.200 73.000 ;
        RECT 63.600 73.000 64.400 73.200 ;
        RECT 72.000 73.000 72.600 74.600 ;
        RECT 63.600 72.400 72.600 73.000 ;
        RECT 72.000 70.600 72.600 72.400 ;
        RECT 73.200 72.000 74.000 79.800 ;
        RECT 83.800 72.600 84.600 79.800 ;
        RECT 88.600 72.600 89.400 79.800 ;
        RECT 90.800 73.800 91.600 79.800 ;
        RECT 91.000 73.200 91.600 73.800 ;
        RECT 94.000 79.200 98.000 79.800 ;
        RECT 94.000 73.800 94.800 79.200 ;
        RECT 95.600 73.800 96.400 78.600 ;
        RECT 97.200 74.000 98.000 79.200 ;
        RECT 99.000 79.200 102.600 79.800 ;
        RECT 99.000 79.000 99.600 79.200 ;
        RECT 94.000 73.200 94.600 73.800 ;
        RECT 91.000 72.600 94.600 73.200 ;
        RECT 95.800 73.400 96.400 73.800 ;
        RECT 98.800 73.400 99.600 79.000 ;
        RECT 102.000 79.000 102.600 79.200 ;
        RECT 95.800 73.000 99.600 73.400 ;
        RECT 100.400 73.000 101.200 78.600 ;
        RECT 102.000 73.000 102.800 79.000 ;
        RECT 95.800 72.800 99.400 73.000 ;
        RECT 73.200 71.200 74.200 72.000 ;
        RECT 82.800 71.800 84.600 72.600 ;
        RECT 87.600 71.800 89.400 72.600 ;
        RECT 100.400 72.400 101.000 73.000 ;
        RECT 103.600 72.400 104.400 79.800 ;
        RECT 100.400 72.200 101.200 72.400 ;
        RECT 42.600 70.000 66.000 70.600 ;
        RECT 72.000 70.000 72.800 70.600 ;
        RECT 42.600 69.800 43.400 70.000 ;
        RECT 44.400 69.600 45.200 70.000 ;
        RECT 47.600 69.600 48.400 70.000 ;
        RECT 54.000 69.600 54.800 70.000 ;
        RECT 65.200 69.400 66.000 70.000 ;
        RECT 41.200 68.200 50.000 69.000 ;
        RECT 50.600 68.600 52.600 69.400 ;
        RECT 56.400 68.600 59.600 69.400 ;
        RECT 41.200 62.200 42.000 68.200 ;
        RECT 43.600 66.800 46.600 67.600 ;
        RECT 45.800 66.200 46.600 66.800 ;
        RECT 51.800 66.200 52.600 68.600 ;
        RECT 54.000 66.800 54.800 68.400 ;
        RECT 59.200 67.800 60.000 68.000 ;
        RECT 55.600 67.200 60.000 67.800 ;
        RECT 55.600 67.000 56.400 67.200 ;
        RECT 62.000 66.400 62.800 69.200 ;
        RECT 67.800 68.600 71.600 69.400 ;
        RECT 67.800 67.400 68.600 68.600 ;
        RECT 72.200 68.000 72.800 70.000 ;
        RECT 55.600 66.200 56.400 66.400 ;
        RECT 45.800 65.400 48.400 66.200 ;
        RECT 51.800 65.600 56.400 66.200 ;
        RECT 61.800 65.600 62.800 66.400 ;
        RECT 66.800 66.800 68.600 67.400 ;
        RECT 71.600 67.400 72.800 68.000 ;
        RECT 66.800 66.200 67.600 66.800 ;
        RECT 47.600 62.200 48.400 65.400 ;
        RECT 65.200 65.400 67.600 66.200 ;
        RECT 49.200 62.200 50.000 65.000 ;
        RECT 50.800 62.200 51.600 65.000 ;
        RECT 52.400 62.200 53.200 65.000 ;
        RECT 55.600 62.200 56.400 65.000 ;
        RECT 58.800 62.200 59.600 65.000 ;
        RECT 60.400 62.200 61.200 65.000 ;
        RECT 62.000 62.200 62.800 65.000 ;
        RECT 63.600 62.200 64.400 65.000 ;
        RECT 65.200 62.200 66.000 65.400 ;
        RECT 71.600 62.200 72.400 67.400 ;
        RECT 73.400 66.800 74.200 71.200 ;
        RECT 83.000 68.400 83.600 71.800 ;
        RECT 84.400 69.600 85.200 71.200 ;
        RECT 87.800 68.400 88.400 71.800 ;
        RECT 97.800 71.600 101.200 72.200 ;
        RECT 103.600 71.800 105.800 72.400 ;
        RECT 89.200 70.300 90.000 71.200 ;
        RECT 95.600 70.300 97.200 70.400 ;
        RECT 89.200 69.700 97.200 70.300 ;
        RECT 89.200 69.600 90.000 69.700 ;
        RECT 95.600 69.600 97.200 69.700 ;
        RECT 74.800 68.300 75.600 68.400 ;
        RECT 82.800 68.300 83.600 68.400 ;
        RECT 74.800 67.700 83.600 68.300 ;
        RECT 74.800 67.600 75.600 67.700 ;
        RECT 82.800 67.600 83.600 67.700 ;
        RECT 87.600 67.600 88.400 68.400 ;
        RECT 94.000 67.600 95.600 68.400 ;
        RECT 73.200 66.000 74.200 66.800 ;
        RECT 73.200 62.200 74.000 66.000 ;
        RECT 81.200 64.800 82.000 66.400 ;
        RECT 83.000 64.200 83.600 67.600 ;
        RECT 86.000 64.800 86.800 66.400 ;
        RECT 87.800 64.400 88.400 67.600 ;
        RECT 92.400 65.600 94.800 66.400 ;
        RECT 97.800 65.000 98.400 71.600 ;
        RECT 105.200 71.200 105.800 71.800 ;
        RECT 105.200 70.400 106.400 71.200 ;
        RECT 103.600 68.800 104.400 70.400 ;
        RECT 105.200 67.400 105.800 70.400 ;
        RECT 94.400 64.400 98.400 65.000 ;
        RECT 82.800 62.200 83.600 64.200 ;
        RECT 87.600 62.200 88.400 64.400 ;
        RECT 94.000 63.600 95.000 64.400 ;
        RECT 97.200 64.200 98.400 64.400 ;
        RECT 103.600 66.800 105.800 67.400 ;
        RECT 94.000 62.200 94.800 63.600 ;
        RECT 97.200 62.200 98.000 64.200 ;
        RECT 103.600 62.200 104.400 66.800 ;
        RECT 1.200 53.800 2.000 59.800 ;
        RECT 7.600 56.600 8.400 59.800 ;
        RECT 9.200 57.000 10.000 59.800 ;
        RECT 10.800 57.000 11.600 59.800 ;
        RECT 12.400 57.000 13.200 59.800 ;
        RECT 15.600 57.000 16.400 59.800 ;
        RECT 18.800 57.000 19.600 59.800 ;
        RECT 20.400 57.000 21.200 59.800 ;
        RECT 22.000 57.000 22.800 59.800 ;
        RECT 23.600 57.000 24.400 59.800 ;
        RECT 5.800 55.800 8.400 56.600 ;
        RECT 25.200 56.600 26.000 59.800 ;
        RECT 11.800 55.800 16.400 56.400 ;
        RECT 5.800 55.200 6.600 55.800 ;
        RECT 3.600 54.400 6.600 55.200 ;
        RECT 1.200 53.000 10.000 53.800 ;
        RECT 11.800 53.400 12.600 55.800 ;
        RECT 15.600 55.600 16.400 55.800 ;
        RECT 21.800 55.600 22.800 56.400 ;
        RECT 25.200 55.800 27.600 56.600 ;
        RECT 14.000 53.600 14.800 55.200 ;
        RECT 15.600 54.800 16.400 55.000 ;
        RECT 15.600 54.200 20.000 54.800 ;
        RECT 19.200 54.000 20.000 54.200 ;
        RECT 1.200 47.400 2.000 53.000 ;
        RECT 10.600 52.600 12.600 53.400 ;
        RECT 16.400 52.600 19.600 53.400 ;
        RECT 22.000 52.800 22.800 55.600 ;
        RECT 26.800 55.200 27.600 55.800 ;
        RECT 26.800 54.600 28.600 55.200 ;
        RECT 27.800 53.400 28.600 54.600 ;
        RECT 31.600 54.600 32.400 59.800 ;
        RECT 33.200 56.000 34.000 59.800 ;
        RECT 33.200 55.200 34.200 56.000 ;
        RECT 41.200 55.800 42.000 59.800 ;
        RECT 45.600 56.200 47.200 59.800 ;
        RECT 41.200 55.200 43.600 55.800 ;
        RECT 31.600 54.000 32.800 54.600 ;
        RECT 27.800 52.600 31.600 53.400 ;
        RECT 2.600 52.000 3.400 52.200 ;
        RECT 4.400 52.000 5.200 52.400 ;
        RECT 7.600 52.000 8.400 52.400 ;
        RECT 25.200 52.000 26.000 52.600 ;
        RECT 32.200 52.000 32.800 54.000 ;
        RECT 2.600 51.400 26.000 52.000 ;
        RECT 32.000 51.400 32.800 52.000 ;
        RECT 33.400 54.300 34.200 55.200 ;
        RECT 42.800 55.000 43.600 55.200 ;
        RECT 44.200 54.800 45.000 55.600 ;
        RECT 44.200 54.400 44.800 54.800 ;
        RECT 41.200 54.300 42.800 54.400 ;
        RECT 33.400 53.700 42.800 54.300 ;
        RECT 32.000 49.600 32.600 51.400 ;
        RECT 33.400 50.800 34.200 53.700 ;
        RECT 41.200 53.600 42.800 53.700 ;
        RECT 44.000 53.600 44.800 54.400 ;
        RECT 45.600 52.800 46.200 56.200 ;
        RECT 50.800 55.800 51.600 59.800 ;
        RECT 52.600 56.400 53.400 57.200 ;
        RECT 46.800 55.400 48.400 55.600 ;
        RECT 46.800 54.800 48.800 55.400 ;
        RECT 49.400 55.200 51.600 55.800 ;
        RECT 52.400 55.600 53.200 56.400 ;
        RECT 54.000 55.800 54.800 59.800 ;
        RECT 49.400 55.000 50.200 55.200 ;
        RECT 48.200 54.400 48.800 54.800 ;
        RECT 46.800 53.400 47.600 54.200 ;
        RECT 48.200 53.800 51.600 54.400 ;
        RECT 50.000 53.600 51.600 53.800 ;
        RECT 45.200 52.400 46.200 52.800 ;
        RECT 34.800 52.300 35.600 52.400 ;
        RECT 44.400 52.300 46.200 52.400 ;
        RECT 34.800 52.200 46.200 52.300 ;
        RECT 47.000 52.800 47.600 53.400 ;
        RECT 47.000 52.200 49.600 52.800 ;
        RECT 34.800 51.700 45.800 52.200 ;
        RECT 48.800 52.000 49.600 52.200 ;
        RECT 52.400 52.200 53.200 52.400 ;
        RECT 54.200 52.200 54.800 55.800 ;
        RECT 60.400 57.800 61.200 59.800 ;
        RECT 60.400 54.400 61.000 57.800 ;
        RECT 62.000 56.300 62.800 57.200 ;
        RECT 64.200 56.400 65.000 59.800 ;
        RECT 70.000 57.800 70.800 59.800 ;
        RECT 64.200 56.300 66.000 56.400 ;
        RECT 62.000 55.700 66.000 56.300 ;
        RECT 62.000 55.600 62.800 55.700 ;
        RECT 55.600 52.800 56.400 54.400 ;
        RECT 60.400 53.600 61.200 54.400 ;
        RECT 57.200 52.200 58.000 52.400 ;
        RECT 34.800 51.600 35.600 51.700 ;
        RECT 44.400 51.600 45.800 51.700 ;
        RECT 52.400 51.600 54.800 52.200 ;
        RECT 56.400 51.600 58.000 52.200 ;
        RECT 10.800 49.400 11.600 49.600 ;
        RECT 6.200 49.000 11.600 49.400 ;
        RECT 5.400 48.800 11.600 49.000 ;
        RECT 12.600 49.000 21.200 49.600 ;
        RECT 2.800 48.000 4.400 48.800 ;
        RECT 5.400 48.200 6.800 48.800 ;
        RECT 12.600 48.200 13.200 49.000 ;
        RECT 20.400 48.800 21.200 49.000 ;
        RECT 23.600 49.000 32.600 49.600 ;
        RECT 23.600 48.800 24.400 49.000 ;
        RECT 3.800 47.600 4.400 48.000 ;
        RECT 7.400 47.600 13.200 48.200 ;
        RECT 13.800 47.600 16.400 48.400 ;
        RECT 1.200 46.800 3.200 47.400 ;
        RECT 3.800 46.800 8.000 47.600 ;
        RECT 2.600 46.200 3.200 46.800 ;
        RECT 2.600 45.600 3.600 46.200 ;
        RECT 2.800 42.200 3.600 45.600 ;
        RECT 6.000 42.200 6.800 46.800 ;
        RECT 9.200 42.200 10.000 45.000 ;
        RECT 10.800 42.200 11.600 45.000 ;
        RECT 12.400 42.200 13.200 47.000 ;
        RECT 15.600 42.200 16.400 47.000 ;
        RECT 18.800 42.200 19.600 48.400 ;
        RECT 26.800 47.600 29.400 48.400 ;
        RECT 22.000 46.800 26.200 47.600 ;
        RECT 20.400 42.200 21.200 45.000 ;
        RECT 22.000 42.200 22.800 45.000 ;
        RECT 23.600 42.200 24.400 45.000 ;
        RECT 26.800 42.200 27.600 47.600 ;
        RECT 32.000 47.400 32.600 49.000 ;
        RECT 30.000 46.800 32.600 47.400 ;
        RECT 33.200 50.000 34.200 50.800 ;
        RECT 45.200 50.200 45.800 51.600 ;
        RECT 46.600 51.400 47.400 51.600 ;
        RECT 46.600 50.800 50.000 51.400 ;
        RECT 49.400 50.200 50.000 50.800 ;
        RECT 52.600 50.200 53.200 51.600 ;
        RECT 56.400 51.200 57.200 51.600 ;
        RECT 58.800 50.800 59.600 52.400 ;
        RECT 60.400 50.200 61.000 53.600 ;
        RECT 30.000 42.200 30.800 46.800 ;
        RECT 33.200 42.200 34.000 50.000 ;
        RECT 41.200 49.600 43.600 50.200 ;
        RECT 45.200 49.600 47.200 50.200 ;
        RECT 41.200 42.200 42.000 49.600 ;
        RECT 42.800 49.400 43.600 49.600 ;
        RECT 45.600 42.200 47.200 49.600 ;
        RECT 49.400 49.600 51.600 50.200 ;
        RECT 49.400 49.400 50.200 49.600 ;
        RECT 50.800 42.200 51.600 49.600 ;
        RECT 52.400 42.200 53.200 50.200 ;
        RECT 54.000 49.600 58.000 50.200 ;
        RECT 54.000 42.200 54.800 49.600 ;
        RECT 57.200 42.200 58.000 49.600 ;
        RECT 59.400 49.400 61.200 50.200 ;
        RECT 59.400 44.400 60.200 49.400 ;
        RECT 63.600 48.800 64.400 50.400 ;
        RECT 58.800 43.600 60.200 44.400 ;
        RECT 59.400 42.200 60.200 43.600 ;
        RECT 65.200 42.200 66.000 55.700 ;
        RECT 68.400 55.600 69.200 57.200 ;
        RECT 66.800 53.600 67.600 55.200 ;
        RECT 70.200 54.400 70.800 57.800 ;
        RECT 73.200 55.600 74.000 57.200 ;
        RECT 74.800 56.300 75.600 59.800 ;
        RECT 82.800 57.800 83.600 59.800 ;
        RECT 81.200 56.300 82.000 56.400 ;
        RECT 74.800 55.700 82.000 56.300 ;
        RECT 70.000 53.600 70.800 54.400 ;
        RECT 70.200 50.200 70.800 53.600 ;
        RECT 71.600 50.800 72.400 52.400 ;
        RECT 70.000 49.400 71.800 50.200 ;
        RECT 71.000 44.400 71.800 49.400 ;
        RECT 70.000 43.600 71.800 44.400 ;
        RECT 71.000 42.200 71.800 43.600 ;
        RECT 74.800 42.200 75.600 55.700 ;
        RECT 81.200 55.600 82.000 55.700 ;
        RECT 82.800 54.400 83.400 57.800 ;
        RECT 84.400 55.600 85.200 57.200 ;
        RECT 76.400 54.300 77.200 54.400 ;
        RECT 82.800 54.300 83.600 54.400 ;
        RECT 76.400 53.700 83.600 54.300 ;
        RECT 87.200 54.200 88.000 59.800 ;
        RECT 92.400 55.200 93.200 59.800 ;
        RECT 97.200 55.200 98.000 59.800 ;
        RECT 102.000 55.200 102.800 59.800 ;
        RECT 92.400 54.600 94.600 55.200 ;
        RECT 97.200 54.600 99.400 55.200 ;
        RECT 102.000 54.600 104.200 55.200 ;
        RECT 76.400 53.600 77.200 53.700 ;
        RECT 82.800 53.600 83.600 53.700 ;
        RECT 86.200 53.800 88.000 54.200 ;
        RECT 86.200 53.600 87.800 53.800 ;
        RECT 81.200 50.800 82.000 52.400 ;
        RECT 82.800 50.200 83.400 53.600 ;
        RECT 86.200 50.400 86.800 53.600 ;
        RECT 88.400 51.600 90.000 52.400 ;
        RECT 92.400 51.600 93.200 53.200 ;
        RECT 94.000 51.600 94.600 54.600 ;
        RECT 97.200 51.600 98.000 53.200 ;
        RECT 98.800 51.600 99.400 54.600 ;
        RECT 102.000 51.600 102.800 53.200 ;
        RECT 103.600 51.600 104.200 54.600 ;
        RECT 81.800 49.400 83.600 50.200 ;
        RECT 86.000 49.600 86.800 50.400 ;
        RECT 90.800 49.600 91.600 51.200 ;
        RECT 94.000 50.800 95.200 51.600 ;
        RECT 98.800 50.800 100.000 51.600 ;
        RECT 103.600 50.800 104.800 51.600 ;
        RECT 94.000 50.200 94.600 50.800 ;
        RECT 98.800 50.200 99.400 50.800 ;
        RECT 103.600 50.200 104.200 50.800 ;
        RECT 92.400 49.600 94.600 50.200 ;
        RECT 97.200 49.600 99.400 50.200 ;
        RECT 102.000 49.600 104.200 50.200 ;
        RECT 81.800 42.200 82.600 49.400 ;
        RECT 86.200 47.000 86.800 49.600 ;
        RECT 87.600 47.600 88.400 49.200 ;
        RECT 86.200 46.400 89.800 47.000 ;
        RECT 86.200 46.200 86.800 46.400 ;
        RECT 86.000 42.200 86.800 46.200 ;
        RECT 89.200 46.200 89.800 46.400 ;
        RECT 89.200 42.200 90.000 46.200 ;
        RECT 92.400 42.200 93.200 49.600 ;
        RECT 97.200 42.200 98.000 49.600 ;
        RECT 102.000 42.200 102.800 49.600 ;
        RECT 2.800 28.300 3.600 39.800 ;
        RECT 7.600 36.400 8.400 39.800 ;
        RECT 7.400 35.800 8.400 36.400 ;
        RECT 7.400 35.200 8.000 35.800 ;
        RECT 10.800 35.200 11.600 39.800 ;
        RECT 14.000 37.000 14.800 39.800 ;
        RECT 15.600 37.000 16.400 39.800 ;
        RECT 6.000 34.600 8.000 35.200 ;
        RECT 6.000 29.000 6.800 34.600 ;
        RECT 8.600 34.400 12.800 35.200 ;
        RECT 17.200 35.000 18.000 39.800 ;
        RECT 20.400 35.000 21.200 39.800 ;
        RECT 8.600 34.000 9.200 34.400 ;
        RECT 7.600 33.200 9.200 34.000 ;
        RECT 12.200 33.800 18.000 34.400 ;
        RECT 10.200 33.200 11.600 33.800 ;
        RECT 10.200 33.000 16.400 33.200 ;
        RECT 11.000 32.600 16.400 33.000 ;
        RECT 15.600 32.400 16.400 32.600 ;
        RECT 17.400 33.000 18.000 33.800 ;
        RECT 18.600 33.600 21.200 34.400 ;
        RECT 23.600 33.600 24.400 39.800 ;
        RECT 25.200 37.000 26.000 39.800 ;
        RECT 26.800 37.000 27.600 39.800 ;
        RECT 28.400 37.000 29.200 39.800 ;
        RECT 26.800 34.400 31.000 35.200 ;
        RECT 31.600 34.400 32.400 39.800 ;
        RECT 34.800 35.200 35.600 39.800 ;
        RECT 34.800 34.600 37.400 35.200 ;
        RECT 31.600 33.600 34.200 34.400 ;
        RECT 25.200 33.000 26.000 33.200 ;
        RECT 17.400 32.400 26.000 33.000 ;
        RECT 28.400 33.000 29.200 33.200 ;
        RECT 36.800 33.000 37.400 34.600 ;
        RECT 28.400 32.400 37.400 33.000 ;
        RECT 36.800 30.600 37.400 32.400 ;
        RECT 38.000 34.300 38.800 39.800 ;
        RECT 41.200 34.300 42.000 34.400 ;
        RECT 38.000 33.700 42.000 34.300 ;
        RECT 38.000 32.000 38.800 33.700 ;
        RECT 41.200 33.600 42.000 33.700 ;
        RECT 46.600 32.600 47.400 39.800 ;
        RECT 52.400 36.400 53.200 39.800 ;
        RECT 52.200 35.800 53.200 36.400 ;
        RECT 52.200 35.200 52.800 35.800 ;
        RECT 55.600 35.200 56.400 39.800 ;
        RECT 58.800 37.000 59.600 39.800 ;
        RECT 60.400 37.000 61.200 39.800 ;
        RECT 50.800 34.600 52.800 35.200 ;
        RECT 38.000 31.200 39.000 32.000 ;
        RECT 46.600 31.800 48.400 32.600 ;
        RECT 7.400 30.000 30.800 30.600 ;
        RECT 36.800 30.000 37.600 30.600 ;
        RECT 7.400 29.800 8.200 30.000 ;
        RECT 9.200 29.600 10.000 30.000 ;
        RECT 12.400 29.600 13.200 30.000 ;
        RECT 30.000 29.400 30.800 30.000 ;
        RECT 4.400 28.300 5.200 28.400 ;
        RECT 2.800 27.700 5.200 28.300 ;
        RECT 2.800 22.200 3.600 27.700 ;
        RECT 4.400 27.600 5.200 27.700 ;
        RECT 6.000 28.200 14.800 29.000 ;
        RECT 15.400 28.600 17.400 29.400 ;
        RECT 21.200 28.600 24.400 29.400 ;
        RECT 6.000 22.200 6.800 28.200 ;
        RECT 8.400 26.800 11.400 27.600 ;
        RECT 10.600 26.200 11.400 26.800 ;
        RECT 16.600 26.200 17.400 28.600 ;
        RECT 18.800 26.800 19.600 28.400 ;
        RECT 24.000 27.800 24.800 28.000 ;
        RECT 20.400 27.200 24.800 27.800 ;
        RECT 20.400 27.000 21.200 27.200 ;
        RECT 26.800 26.400 27.600 29.200 ;
        RECT 32.600 28.600 36.400 29.400 ;
        RECT 32.600 27.400 33.400 28.600 ;
        RECT 37.000 28.000 37.600 30.000 ;
        RECT 20.400 26.200 21.200 26.400 ;
        RECT 10.600 25.400 13.200 26.200 ;
        RECT 16.600 25.600 21.200 26.200 ;
        RECT 26.600 25.600 27.600 26.400 ;
        RECT 31.600 26.800 33.400 27.400 ;
        RECT 36.400 27.400 37.600 28.000 ;
        RECT 31.600 26.200 32.400 26.800 ;
        RECT 12.400 22.200 13.200 25.400 ;
        RECT 30.000 25.400 32.400 26.200 ;
        RECT 14.000 22.200 14.800 25.000 ;
        RECT 15.600 22.200 16.400 25.000 ;
        RECT 17.200 22.200 18.000 25.000 ;
        RECT 20.400 22.200 21.200 25.000 ;
        RECT 23.600 22.200 24.400 25.000 ;
        RECT 25.200 22.200 26.000 25.000 ;
        RECT 26.800 22.200 27.600 25.000 ;
        RECT 28.400 22.200 29.200 25.000 ;
        RECT 30.000 22.200 30.800 25.400 ;
        RECT 36.400 22.200 37.200 27.400 ;
        RECT 38.200 26.800 39.000 31.200 ;
        RECT 46.000 29.600 46.800 31.200 ;
        RECT 47.600 28.400 48.200 31.800 ;
        RECT 50.800 29.000 51.600 34.600 ;
        RECT 53.400 34.400 57.600 35.200 ;
        RECT 62.000 35.000 62.800 39.800 ;
        RECT 65.200 35.000 66.000 39.800 ;
        RECT 53.400 34.000 54.000 34.400 ;
        RECT 52.400 33.200 54.000 34.000 ;
        RECT 57.000 33.800 62.800 34.400 ;
        RECT 55.000 33.200 56.400 33.800 ;
        RECT 55.000 33.000 61.200 33.200 ;
        RECT 55.800 32.600 61.200 33.000 ;
        RECT 60.400 32.400 61.200 32.600 ;
        RECT 62.200 33.000 62.800 33.800 ;
        RECT 63.400 33.600 66.000 34.400 ;
        RECT 68.400 33.600 69.200 39.800 ;
        RECT 70.000 37.000 70.800 39.800 ;
        RECT 71.600 37.000 72.400 39.800 ;
        RECT 73.200 37.000 74.000 39.800 ;
        RECT 71.600 34.400 75.800 35.200 ;
        RECT 76.400 34.400 77.200 39.800 ;
        RECT 79.600 35.200 80.400 39.800 ;
        RECT 79.600 34.600 82.200 35.200 ;
        RECT 76.400 33.600 79.000 34.400 ;
        RECT 70.000 33.000 70.800 33.200 ;
        RECT 62.200 32.400 70.800 33.000 ;
        RECT 73.200 33.000 74.000 33.200 ;
        RECT 81.600 33.000 82.200 34.600 ;
        RECT 73.200 32.400 82.200 33.000 ;
        RECT 81.600 30.600 82.200 32.400 ;
        RECT 82.800 34.300 83.600 39.800 ;
        RECT 90.800 35.800 91.600 39.800 ;
        RECT 91.000 35.600 91.600 35.800 ;
        RECT 94.000 35.800 94.800 39.800 ;
        RECT 94.000 35.600 94.600 35.800 ;
        RECT 91.000 35.000 94.600 35.600 ;
        RECT 84.400 34.300 85.200 34.400 ;
        RECT 82.800 33.700 85.200 34.300 ;
        RECT 82.800 32.000 83.600 33.700 ;
        RECT 84.400 33.600 85.200 33.700 ;
        RECT 91.000 32.400 91.600 35.000 ;
        RECT 92.400 32.800 93.200 34.400 ;
        RECT 82.800 31.200 83.800 32.000 ;
        RECT 90.800 31.600 91.600 32.400 ;
        RECT 52.200 30.000 75.600 30.600 ;
        RECT 81.600 30.000 82.400 30.600 ;
        RECT 52.200 29.800 53.000 30.000 ;
        RECT 54.000 29.600 54.800 30.000 ;
        RECT 55.600 29.600 56.400 30.000 ;
        RECT 57.200 29.600 58.000 30.000 ;
        RECT 74.800 29.400 75.600 30.000 ;
        RECT 39.600 28.300 40.400 28.400 ;
        RECT 47.600 28.300 48.400 28.400 ;
        RECT 39.600 27.700 48.400 28.300 ;
        RECT 39.600 27.600 40.400 27.700 ;
        RECT 47.600 27.600 48.400 27.700 ;
        RECT 50.800 28.200 59.600 29.000 ;
        RECT 60.200 28.600 62.200 29.400 ;
        RECT 66.000 28.600 69.200 29.400 ;
        RECT 38.000 26.000 39.000 26.800 ;
        RECT 38.000 22.200 38.800 26.000 ;
        RECT 47.600 24.200 48.200 27.600 ;
        RECT 49.200 24.800 50.000 26.400 ;
        RECT 47.600 22.200 48.400 24.200 ;
        RECT 50.800 22.200 51.600 28.200 ;
        RECT 53.200 26.800 56.200 27.600 ;
        RECT 55.400 26.200 56.200 26.800 ;
        RECT 61.400 26.200 62.200 28.600 ;
        RECT 63.600 26.800 64.400 28.400 ;
        RECT 68.800 27.800 69.600 28.000 ;
        RECT 65.200 27.200 69.600 27.800 ;
        RECT 65.200 27.000 66.000 27.200 ;
        RECT 71.600 26.400 72.400 29.200 ;
        RECT 77.400 28.600 81.200 29.400 ;
        RECT 77.400 27.400 78.200 28.600 ;
        RECT 81.800 28.000 82.400 30.000 ;
        RECT 65.200 26.200 66.000 26.400 ;
        RECT 55.400 25.400 58.000 26.200 ;
        RECT 61.400 25.600 66.000 26.200 ;
        RECT 71.400 25.600 72.400 26.400 ;
        RECT 76.400 26.800 78.200 27.400 ;
        RECT 81.200 27.400 82.400 28.000 ;
        RECT 76.400 26.200 77.200 26.800 ;
        RECT 57.200 22.200 58.000 25.400 ;
        RECT 74.800 25.400 77.200 26.200 ;
        RECT 58.800 22.200 59.600 25.000 ;
        RECT 60.400 22.200 61.200 25.000 ;
        RECT 62.000 22.200 62.800 25.000 ;
        RECT 65.200 22.200 66.000 25.000 ;
        RECT 68.400 22.200 69.200 25.000 ;
        RECT 70.000 22.200 70.800 25.000 ;
        RECT 71.600 22.200 72.400 25.000 ;
        RECT 73.200 22.200 74.000 25.000 ;
        RECT 74.800 22.200 75.600 25.400 ;
        RECT 81.200 22.200 82.000 27.400 ;
        RECT 83.000 26.800 83.800 31.200 ;
        RECT 91.000 28.400 91.600 31.600 ;
        RECT 95.600 30.800 96.400 32.400 ;
        RECT 93.200 29.600 94.800 30.400 ;
        RECT 91.000 28.200 92.600 28.400 ;
        RECT 91.000 27.800 92.800 28.200 ;
        RECT 82.800 26.300 83.800 26.800 ;
        RECT 89.200 26.300 90.000 26.400 ;
        RECT 82.800 25.700 90.000 26.300 ;
        RECT 82.800 22.200 83.600 25.700 ;
        RECT 89.200 25.600 90.000 25.700 ;
        RECT 92.000 24.400 92.800 27.800 ;
        RECT 92.000 23.600 93.200 24.400 ;
        RECT 92.000 22.200 92.800 23.600 ;
        RECT 97.200 22.200 98.000 39.800 ;
        RECT 100.400 32.400 101.200 39.800 ;
        RECT 105.200 32.400 106.000 39.800 ;
        RECT 100.400 31.800 102.600 32.400 ;
        RECT 105.200 31.800 107.400 32.400 ;
        RECT 102.000 31.200 102.600 31.800 ;
        RECT 106.800 31.200 107.400 31.800 ;
        RECT 102.000 30.400 103.200 31.200 ;
        RECT 106.800 30.400 108.000 31.200 ;
        RECT 100.400 28.800 101.200 30.400 ;
        RECT 102.000 27.400 102.600 30.400 ;
        RECT 105.200 28.800 106.000 30.400 ;
        RECT 106.800 27.400 107.400 30.400 ;
        RECT 100.400 26.800 102.600 27.400 ;
        RECT 105.200 26.800 107.400 27.400 ;
        RECT 98.800 24.800 99.600 26.400 ;
        RECT 100.400 22.200 101.200 26.800 ;
        RECT 105.200 22.200 106.000 26.800 ;
        RECT 1.200 13.800 2.000 19.800 ;
        RECT 7.600 16.600 8.400 19.800 ;
        RECT 9.200 17.000 10.000 19.800 ;
        RECT 10.800 17.000 11.600 19.800 ;
        RECT 12.400 17.000 13.200 19.800 ;
        RECT 15.600 17.000 16.400 19.800 ;
        RECT 18.800 17.000 19.600 19.800 ;
        RECT 20.400 17.000 21.200 19.800 ;
        RECT 22.000 17.000 22.800 19.800 ;
        RECT 23.600 17.000 24.400 19.800 ;
        RECT 5.800 15.800 8.400 16.600 ;
        RECT 25.200 16.600 26.000 19.800 ;
        RECT 11.800 15.800 16.400 16.400 ;
        RECT 5.800 15.200 6.600 15.800 ;
        RECT 3.600 14.400 6.600 15.200 ;
        RECT 1.200 13.000 10.000 13.800 ;
        RECT 11.800 13.400 12.600 15.800 ;
        RECT 15.600 15.600 16.400 15.800 ;
        RECT 21.800 15.600 22.800 16.400 ;
        RECT 25.200 15.800 27.600 16.600 ;
        RECT 14.000 13.600 14.800 15.200 ;
        RECT 15.600 14.800 16.400 15.000 ;
        RECT 15.600 14.200 20.000 14.800 ;
        RECT 19.200 14.000 20.000 14.200 ;
        RECT 1.200 7.400 2.000 13.000 ;
        RECT 10.600 12.600 12.600 13.400 ;
        RECT 16.400 12.600 19.600 13.400 ;
        RECT 22.000 12.800 22.800 15.600 ;
        RECT 26.800 15.200 27.600 15.800 ;
        RECT 26.800 14.600 28.600 15.200 ;
        RECT 27.800 13.400 28.600 14.600 ;
        RECT 31.600 14.600 32.400 19.800 ;
        RECT 33.200 16.000 34.000 19.800 ;
        RECT 33.200 15.200 34.200 16.000 ;
        RECT 41.200 15.800 42.000 19.800 ;
        RECT 45.600 16.200 47.200 19.800 ;
        RECT 41.200 15.200 43.600 15.800 ;
        RECT 31.600 14.000 32.800 14.600 ;
        RECT 27.800 12.600 31.600 13.400 ;
        RECT 2.600 12.000 3.400 12.200 ;
        RECT 4.400 12.000 5.200 12.400 ;
        RECT 7.600 12.000 8.400 12.400 ;
        RECT 25.200 12.000 26.000 12.600 ;
        RECT 32.200 12.000 32.800 14.000 ;
        RECT 2.600 11.400 26.000 12.000 ;
        RECT 32.000 11.400 32.800 12.000 ;
        RECT 33.400 14.300 34.200 15.200 ;
        RECT 42.800 15.000 43.600 15.200 ;
        RECT 44.200 14.800 45.000 15.600 ;
        RECT 44.200 14.400 44.800 14.800 ;
        RECT 41.200 14.300 42.800 14.400 ;
        RECT 33.400 13.700 42.800 14.300 ;
        RECT 32.000 9.600 32.600 11.400 ;
        RECT 33.400 10.800 34.200 13.700 ;
        RECT 41.200 13.600 42.800 13.700 ;
        RECT 44.000 13.600 44.800 14.400 ;
        RECT 45.600 12.800 46.200 16.200 ;
        RECT 50.800 15.800 51.600 19.800 ;
        RECT 46.800 15.400 48.400 15.600 ;
        RECT 46.800 14.800 48.800 15.400 ;
        RECT 49.400 15.200 51.600 15.800 ;
        RECT 49.400 15.000 50.200 15.200 ;
        RECT 48.200 14.400 48.800 14.800 ;
        RECT 46.800 13.400 47.600 14.200 ;
        RECT 48.200 13.800 51.600 14.400 ;
        RECT 50.000 13.600 51.600 13.800 ;
        RECT 52.400 13.800 53.200 19.800 ;
        RECT 58.800 16.600 59.600 19.800 ;
        RECT 60.400 17.000 61.200 19.800 ;
        RECT 62.000 17.000 62.800 19.800 ;
        RECT 63.600 17.000 64.400 19.800 ;
        RECT 66.800 17.000 67.600 19.800 ;
        RECT 70.000 17.000 70.800 19.800 ;
        RECT 71.600 17.000 72.400 19.800 ;
        RECT 73.200 17.000 74.000 19.800 ;
        RECT 74.800 17.000 75.600 19.800 ;
        RECT 57.000 15.800 59.600 16.600 ;
        RECT 76.400 16.600 77.200 19.800 ;
        RECT 63.000 15.800 67.600 16.400 ;
        RECT 57.000 15.200 57.800 15.800 ;
        RECT 54.800 14.400 57.800 15.200 ;
        RECT 45.200 12.400 46.200 12.800 ;
        RECT 34.800 12.300 35.600 12.400 ;
        RECT 44.400 12.300 46.200 12.400 ;
        RECT 34.800 12.200 46.200 12.300 ;
        RECT 47.000 12.800 47.600 13.400 ;
        RECT 52.400 13.000 61.200 13.800 ;
        RECT 63.000 13.400 63.800 15.800 ;
        RECT 66.800 15.600 67.600 15.800 ;
        RECT 73.000 15.600 74.000 16.400 ;
        RECT 76.400 15.800 78.800 16.600 ;
        RECT 65.200 13.600 66.000 15.200 ;
        RECT 66.800 14.800 67.600 15.000 ;
        RECT 66.800 14.200 71.200 14.800 ;
        RECT 70.400 14.000 71.200 14.200 ;
        RECT 47.000 12.200 49.600 12.800 ;
        RECT 34.800 11.700 45.800 12.200 ;
        RECT 48.800 12.000 49.600 12.200 ;
        RECT 34.800 11.600 35.600 11.700 ;
        RECT 44.400 11.600 45.800 11.700 ;
        RECT 10.800 9.400 11.600 9.600 ;
        RECT 6.200 9.000 11.600 9.400 ;
        RECT 5.400 8.800 11.600 9.000 ;
        RECT 12.600 9.000 21.200 9.600 ;
        RECT 2.800 8.000 4.400 8.800 ;
        RECT 5.400 8.200 6.800 8.800 ;
        RECT 12.600 8.200 13.200 9.000 ;
        RECT 20.400 8.800 21.200 9.000 ;
        RECT 23.600 9.000 32.600 9.600 ;
        RECT 23.600 8.800 24.400 9.000 ;
        RECT 3.800 7.600 4.400 8.000 ;
        RECT 7.400 7.600 13.200 8.200 ;
        RECT 13.800 7.600 16.400 8.400 ;
        RECT 1.200 6.800 3.200 7.400 ;
        RECT 3.800 6.800 8.000 7.600 ;
        RECT 2.600 6.200 3.200 6.800 ;
        RECT 2.600 5.600 3.600 6.200 ;
        RECT 2.800 2.200 3.600 5.600 ;
        RECT 6.000 2.200 6.800 6.800 ;
        RECT 9.200 2.200 10.000 5.000 ;
        RECT 10.800 2.200 11.600 5.000 ;
        RECT 12.400 2.200 13.200 7.000 ;
        RECT 15.600 2.200 16.400 7.000 ;
        RECT 18.800 2.200 19.600 8.400 ;
        RECT 26.800 7.600 29.400 8.400 ;
        RECT 22.000 6.800 26.200 7.600 ;
        RECT 20.400 2.200 21.200 5.000 ;
        RECT 22.000 2.200 22.800 5.000 ;
        RECT 23.600 2.200 24.400 5.000 ;
        RECT 26.800 2.200 27.600 7.600 ;
        RECT 32.000 7.400 32.600 9.000 ;
        RECT 30.000 6.800 32.600 7.400 ;
        RECT 33.200 10.000 34.200 10.800 ;
        RECT 45.200 10.200 45.800 11.600 ;
        RECT 46.600 11.400 47.400 11.600 ;
        RECT 46.600 10.800 50.000 11.400 ;
        RECT 49.400 10.200 50.000 10.800 ;
        RECT 30.000 2.200 30.800 6.800 ;
        RECT 33.200 2.200 34.000 10.000 ;
        RECT 41.200 9.600 43.600 10.200 ;
        RECT 45.200 9.600 47.200 10.200 ;
        RECT 41.200 2.200 42.000 9.600 ;
        RECT 42.800 9.400 43.600 9.600 ;
        RECT 45.600 2.200 47.200 9.600 ;
        RECT 49.400 9.600 51.600 10.200 ;
        RECT 49.400 9.400 50.200 9.600 ;
        RECT 50.800 2.200 51.600 9.600 ;
        RECT 52.400 7.400 53.200 13.000 ;
        RECT 61.800 12.600 63.800 13.400 ;
        RECT 67.600 12.600 70.800 13.400 ;
        RECT 73.200 12.800 74.000 15.600 ;
        RECT 78.000 15.200 78.800 15.800 ;
        RECT 78.000 14.600 79.800 15.200 ;
        RECT 79.000 13.400 79.800 14.600 ;
        RECT 82.800 14.600 83.600 19.800 ;
        RECT 84.400 16.300 85.200 19.800 ;
        RECT 86.000 16.300 86.800 16.400 ;
        RECT 84.400 15.700 86.800 16.300 ;
        RECT 84.400 15.200 85.400 15.700 ;
        RECT 86.000 15.600 86.800 15.700 ;
        RECT 89.200 16.300 90.000 16.400 ;
        RECT 92.400 16.300 93.200 17.200 ;
        RECT 89.200 15.700 93.200 16.300 ;
        RECT 89.200 15.600 90.000 15.700 ;
        RECT 92.400 15.600 93.200 15.700 ;
        RECT 82.800 14.000 84.000 14.600 ;
        RECT 79.000 12.600 82.800 13.400 ;
        RECT 53.800 12.000 54.600 12.200 ;
        RECT 55.600 12.000 56.400 12.400 ;
        RECT 58.800 12.000 59.600 12.400 ;
        RECT 76.400 12.000 77.200 12.600 ;
        RECT 83.400 12.000 84.000 14.000 ;
        RECT 53.800 11.400 77.200 12.000 ;
        RECT 83.200 11.400 84.000 12.000 ;
        RECT 83.200 9.600 83.800 11.400 ;
        RECT 84.600 10.800 85.400 15.200 ;
        RECT 62.000 9.400 62.800 9.600 ;
        RECT 57.400 9.000 62.800 9.400 ;
        RECT 56.600 8.800 62.800 9.000 ;
        RECT 63.800 9.000 72.400 9.600 ;
        RECT 54.000 8.000 55.600 8.800 ;
        RECT 56.600 8.200 58.000 8.800 ;
        RECT 63.800 8.200 64.400 9.000 ;
        RECT 71.600 8.800 72.400 9.000 ;
        RECT 74.800 9.000 83.800 9.600 ;
        RECT 74.800 8.800 75.600 9.000 ;
        RECT 55.000 7.600 55.600 8.000 ;
        RECT 58.600 7.600 64.400 8.200 ;
        RECT 65.000 7.600 67.600 8.400 ;
        RECT 52.400 6.800 54.400 7.400 ;
        RECT 55.000 6.800 59.200 7.600 ;
        RECT 53.800 6.200 54.400 6.800 ;
        RECT 53.800 5.600 54.800 6.200 ;
        RECT 54.000 2.200 54.800 5.600 ;
        RECT 57.200 2.200 58.000 6.800 ;
        RECT 60.400 2.200 61.200 5.000 ;
        RECT 62.000 2.200 62.800 5.000 ;
        RECT 63.600 2.200 64.400 7.000 ;
        RECT 66.800 2.200 67.600 7.000 ;
        RECT 70.000 2.200 70.800 8.400 ;
        RECT 78.000 7.600 80.600 8.400 ;
        RECT 73.200 6.800 77.400 7.600 ;
        RECT 71.600 2.200 72.400 5.000 ;
        RECT 73.200 2.200 74.000 5.000 ;
        RECT 74.800 2.200 75.600 5.000 ;
        RECT 78.000 2.200 78.800 7.600 ;
        RECT 83.200 7.400 83.800 9.000 ;
        RECT 81.200 6.800 83.800 7.400 ;
        RECT 84.400 10.000 85.400 10.800 ;
        RECT 81.200 2.200 82.000 6.800 ;
        RECT 84.400 2.200 85.200 10.000 ;
        RECT 94.000 2.200 94.800 19.800 ;
        RECT 96.200 16.400 97.000 19.800 ;
        RECT 96.200 15.800 98.000 16.400 ;
        RECT 95.600 14.300 96.400 14.400 ;
        RECT 97.200 14.300 98.000 15.800 ;
        RECT 100.400 15.600 101.200 17.200 ;
        RECT 95.600 13.700 98.000 14.300 ;
        RECT 95.600 13.600 96.400 13.700 ;
        RECT 95.600 8.800 96.400 10.400 ;
        RECT 97.200 2.200 98.000 13.700 ;
        RECT 98.800 13.600 99.600 15.200 ;
        RECT 102.000 14.300 102.800 19.800 ;
        RECT 103.600 16.000 104.400 19.800 ;
        RECT 106.800 16.000 107.600 19.800 ;
        RECT 103.600 15.800 107.600 16.000 ;
        RECT 108.400 15.800 109.200 19.800 ;
        RECT 103.800 15.400 107.400 15.800 ;
        RECT 104.400 14.400 105.200 14.800 ;
        RECT 108.400 14.400 109.000 15.800 ;
        RECT 103.600 14.300 105.200 14.400 ;
        RECT 102.000 13.800 105.200 14.300 ;
        RECT 102.000 13.700 104.400 13.800 ;
        RECT 102.000 2.200 102.800 13.700 ;
        RECT 103.600 13.600 104.400 13.700 ;
        RECT 106.600 13.600 109.200 14.400 ;
        RECT 103.600 12.300 104.400 12.400 ;
        RECT 105.200 12.300 106.000 13.200 ;
        RECT 103.600 11.700 106.000 12.300 ;
        RECT 103.600 11.600 104.400 11.700 ;
        RECT 105.200 11.600 106.000 11.700 ;
        RECT 106.600 10.200 107.200 13.600 ;
        RECT 108.400 10.200 109.200 10.400 ;
        RECT 106.200 9.600 107.200 10.200 ;
        RECT 107.800 9.600 109.200 10.200 ;
        RECT 106.200 2.200 107.000 9.600 ;
        RECT 107.800 8.400 108.400 9.600 ;
        RECT 107.600 7.600 108.400 8.400 ;
      LAYER via1 ;
        RECT 7.600 91.600 8.400 92.400 ;
        RECT 20.400 95.600 21.200 96.400 ;
        RECT 15.600 91.600 16.400 92.400 ;
        RECT 15.600 83.600 16.400 84.400 ;
        RECT 39.600 93.000 40.400 93.800 ;
        RECT 49.200 92.600 50.000 93.400 ;
        RECT 55.600 91.600 56.400 92.400 ;
        RECT 73.200 94.800 74.000 95.600 ;
        RECT 76.400 93.600 77.200 94.400 ;
        RECT 86.000 93.600 86.800 94.400 ;
        RECT 41.200 88.800 42.000 89.600 ;
        RECT 46.000 87.600 46.800 88.400 ;
        RECT 42.800 86.200 43.600 87.000 ;
        RECT 39.600 84.200 40.400 85.000 ;
        RECT 41.200 84.200 42.000 85.000 ;
        RECT 46.000 86.200 46.800 87.000 ;
        RECT 49.200 86.200 50.000 87.000 ;
        RECT 50.800 84.200 51.600 85.000 ;
        RECT 52.400 84.200 53.200 85.000 ;
        RECT 54.000 84.200 54.800 85.000 ;
        RECT 87.600 91.600 88.400 92.400 ;
        RECT 100.400 93.600 101.200 94.400 ;
        RECT 95.600 87.600 96.400 88.400 ;
        RECT 94.000 83.600 94.800 84.400 ;
        RECT 102.000 89.600 102.800 90.400 ;
        RECT 103.600 83.600 104.400 84.400 ;
        RECT 2.800 77.600 3.600 78.400 ;
        RECT 14.000 74.400 14.800 75.200 ;
        RECT 17.200 75.000 18.000 75.800 ;
        RECT 12.400 72.400 13.200 73.200 ;
        RECT 10.800 69.600 11.600 70.400 ;
        RECT 22.000 67.600 22.800 68.400 ;
        RECT 12.400 64.200 13.200 65.000 ;
        RECT 14.000 64.200 14.800 65.000 ;
        RECT 15.600 64.200 16.400 65.000 ;
        RECT 17.200 64.200 18.000 65.000 ;
        RECT 20.400 64.200 21.200 65.000 ;
        RECT 23.600 64.200 24.400 65.000 ;
        RECT 25.200 64.200 26.000 65.000 ;
        RECT 26.800 64.200 27.600 65.000 ;
        RECT 58.800 75.000 59.600 75.800 ;
        RECT 55.600 73.600 56.400 74.400 ;
        RECT 73.200 77.600 74.000 78.400 ;
        RECT 60.400 72.400 61.200 73.200 ;
        RECT 49.200 68.200 50.000 69.000 ;
        RECT 58.800 68.600 59.600 69.400 ;
        RECT 54.000 67.600 54.800 68.400 ;
        RECT 49.200 64.200 50.000 65.000 ;
        RECT 50.800 64.200 51.600 65.000 ;
        RECT 52.400 64.200 53.200 65.000 ;
        RECT 55.600 64.200 56.400 65.000 ;
        RECT 58.800 64.200 59.600 65.000 ;
        RECT 60.400 64.200 61.200 65.000 ;
        RECT 62.000 64.200 62.800 65.000 ;
        RECT 63.600 64.200 64.400 65.000 ;
        RECT 81.200 65.600 82.000 66.400 ;
        RECT 86.000 65.600 86.800 66.400 ;
        RECT 94.000 65.600 94.800 66.400 ;
        RECT 103.600 69.600 104.400 70.400 ;
        RECT 87.600 63.600 88.400 64.400 ;
        RECT 9.200 53.000 10.000 53.800 ;
        RECT 18.800 52.600 19.600 53.400 ;
        RECT 4.400 51.600 5.200 52.400 ;
        RECT 47.600 54.800 48.400 55.600 ;
        RECT 50.800 53.600 51.600 54.400 ;
        RECT 65.200 55.600 66.000 56.400 ;
        RECT 55.600 53.600 56.400 54.400 ;
        RECT 10.800 48.800 11.600 49.600 ;
        RECT 15.600 47.600 16.400 48.400 ;
        RECT 12.400 46.200 13.200 47.000 ;
        RECT 9.200 44.200 10.000 45.000 ;
        RECT 10.800 44.200 11.600 45.000 ;
        RECT 15.600 46.200 16.400 47.000 ;
        RECT 18.800 46.200 19.600 47.000 ;
        RECT 20.400 44.200 21.200 45.000 ;
        RECT 22.000 44.200 22.800 45.000 ;
        RECT 23.600 44.200 24.400 45.000 ;
        RECT 57.200 51.600 58.000 52.400 ;
        RECT 58.800 51.600 59.600 52.400 ;
        RECT 52.400 43.600 53.200 44.400 ;
        RECT 63.600 49.600 64.400 50.400 ;
        RECT 71.600 51.600 72.400 52.400 ;
        RECT 81.200 51.600 82.000 52.400 ;
        RECT 89.200 51.600 90.000 52.400 ;
        RECT 89.200 43.600 90.000 44.400 ;
        RECT 23.600 35.000 24.400 35.800 ;
        RECT 20.400 33.600 21.200 34.400 ;
        RECT 25.200 32.400 26.000 33.200 ;
        RECT 30.000 29.600 30.800 30.400 ;
        RECT 14.000 28.200 14.800 29.000 ;
        RECT 23.600 28.600 24.400 29.400 ;
        RECT 18.800 27.600 19.600 28.400 ;
        RECT 14.000 24.200 14.800 25.000 ;
        RECT 15.600 24.200 16.400 25.000 ;
        RECT 17.200 24.200 18.000 25.000 ;
        RECT 20.400 24.200 21.200 25.000 ;
        RECT 23.600 24.200 24.400 25.000 ;
        RECT 25.200 24.200 26.000 25.000 ;
        RECT 26.800 24.200 27.600 25.000 ;
        RECT 28.400 24.200 29.200 25.000 ;
        RECT 68.400 35.000 69.200 35.800 ;
        RECT 65.200 33.600 66.000 34.400 ;
        RECT 70.000 32.400 70.800 33.200 ;
        RECT 92.400 33.600 93.200 34.400 ;
        RECT 58.800 28.200 59.600 29.000 ;
        RECT 68.400 28.600 69.200 29.400 ;
        RECT 49.200 25.600 50.000 26.400 ;
        RECT 63.600 27.600 64.400 28.400 ;
        RECT 58.800 24.200 59.600 25.000 ;
        RECT 60.400 24.200 61.200 25.000 ;
        RECT 62.000 24.200 62.800 25.000 ;
        RECT 65.200 24.200 66.000 25.000 ;
        RECT 68.400 24.200 69.200 25.000 ;
        RECT 70.000 24.200 70.800 25.000 ;
        RECT 71.600 24.200 72.400 25.000 ;
        RECT 73.200 24.200 74.000 25.000 ;
        RECT 95.600 31.600 96.400 32.400 ;
        RECT 94.000 29.600 94.800 30.400 ;
        RECT 97.200 29.600 98.000 30.400 ;
        RECT 92.400 23.600 93.200 24.400 ;
        RECT 100.400 29.600 101.200 30.400 ;
        RECT 105.200 29.600 106.000 30.400 ;
        RECT 98.800 25.600 99.600 26.400 ;
        RECT 9.200 13.000 10.000 13.800 ;
        RECT 18.800 12.600 19.600 13.400 ;
        RECT 4.400 11.600 5.200 12.400 ;
        RECT 47.600 14.800 48.400 15.600 ;
        RECT 50.800 13.600 51.600 14.400 ;
        RECT 60.400 13.000 61.200 13.800 ;
        RECT 10.800 8.800 11.600 9.600 ;
        RECT 15.600 7.600 16.400 8.400 ;
        RECT 12.400 6.200 13.200 7.000 ;
        RECT 9.200 4.200 10.000 5.000 ;
        RECT 10.800 4.200 11.600 5.000 ;
        RECT 15.600 6.200 16.400 7.000 ;
        RECT 18.800 6.200 19.600 7.000 ;
        RECT 20.400 4.200 21.200 5.000 ;
        RECT 22.000 4.200 22.800 5.000 ;
        RECT 23.600 4.200 24.400 5.000 ;
        RECT 70.000 12.600 70.800 13.400 ;
        RECT 94.000 17.600 94.800 18.400 ;
        RECT 55.600 11.600 56.400 12.400 ;
        RECT 62.000 8.800 62.800 9.600 ;
        RECT 66.800 7.600 67.600 8.400 ;
        RECT 63.600 6.200 64.400 7.000 ;
        RECT 60.400 4.200 61.200 5.000 ;
        RECT 62.000 4.200 62.800 5.000 ;
        RECT 66.800 6.200 67.600 7.000 ;
        RECT 70.000 6.200 70.800 7.000 ;
        RECT 71.600 4.200 72.400 5.000 ;
        RECT 73.200 4.200 74.000 5.000 ;
        RECT 74.800 4.200 75.600 5.000 ;
        RECT 95.600 9.600 96.400 10.400 ;
        RECT 106.800 13.600 107.600 14.400 ;
        RECT 108.400 9.600 109.200 10.400 ;
      LAYER metal2 ;
        RECT 20.400 95.600 21.200 96.400 ;
        RECT 6.000 93.600 6.800 94.400 ;
        RECT 15.600 93.600 16.400 94.400 ;
        RECT 6.100 92.400 6.700 93.600 ;
        RECT 15.700 92.400 16.300 93.600 ;
        RECT 2.800 91.600 3.600 92.400 ;
        RECT 6.000 91.600 6.800 92.400 ;
        RECT 7.600 91.600 8.400 92.400 ;
        RECT 15.600 91.600 16.400 92.400 ;
        RECT 22.000 91.600 22.800 92.400 ;
        RECT 2.900 78.400 3.500 91.600 ;
        RECT 15.600 83.600 16.400 84.400 ;
        RECT 39.600 84.200 40.400 97.800 ;
        RECT 41.200 84.200 42.000 97.800 ;
        RECT 42.800 86.200 43.600 97.800 ;
        RECT 44.400 93.600 45.200 94.400 ;
        RECT 44.500 92.400 45.100 93.600 ;
        RECT 44.400 91.600 45.200 92.400 ;
        RECT 46.000 86.200 46.800 97.800 ;
        RECT 49.200 86.200 50.000 97.800 ;
        RECT 50.800 84.200 51.600 97.800 ;
        RECT 52.400 84.200 53.200 97.800 ;
        RECT 54.000 84.200 54.800 97.800 ;
        RECT 68.400 95.000 69.200 95.800 ;
        RECT 69.800 95.000 74.000 95.600 ;
        RECT 75.000 95.000 75.800 95.800 ;
        RECT 76.400 95.600 77.200 96.400 ;
        RECT 82.800 95.600 83.600 96.400 ;
        RECT 98.800 95.600 99.600 96.400 ;
        RECT 102.000 95.600 102.800 96.400 ;
        RECT 106.800 95.600 107.600 96.400 ;
        RECT 66.800 93.600 67.600 94.400 ;
        RECT 68.400 94.200 69.000 95.000 ;
        RECT 69.800 94.800 70.600 95.000 ;
        RECT 73.200 94.800 74.000 95.000 ;
        RECT 68.400 93.600 73.200 94.200 ;
        RECT 66.900 92.400 67.500 93.600 ;
        RECT 55.600 91.600 56.400 92.400 ;
        RECT 65.200 91.600 66.000 92.400 ;
        RECT 66.800 91.600 67.600 92.400 ;
        RECT 15.700 80.400 16.300 83.600 ;
        RECT 55.700 82.300 56.300 91.600 ;
        RECT 68.400 90.200 69.000 93.600 ;
        RECT 72.400 93.400 73.200 93.600 ;
        RECT 75.200 90.200 75.800 95.000 ;
        RECT 76.500 94.400 77.100 95.600 ;
        RECT 76.400 93.600 77.200 94.400 ;
        RECT 68.400 89.400 69.200 90.200 ;
        RECT 75.000 89.400 75.800 90.200 ;
        RECT 54.100 81.700 56.300 82.300 ;
        RECT 15.600 79.600 16.400 80.400 ;
        RECT 22.000 79.600 22.800 80.400 ;
        RECT 2.800 77.600 3.600 78.400 ;
        RECT 4.400 69.600 5.200 70.400 ;
        RECT 10.800 69.600 11.600 70.400 ;
        RECT 4.500 52.400 5.100 69.600 ;
        RECT 12.400 64.200 13.200 77.800 ;
        RECT 14.000 64.200 14.800 77.800 ;
        RECT 15.600 64.200 16.400 77.800 ;
        RECT 17.200 64.200 18.000 75.800 ;
        RECT 20.400 64.200 21.200 75.800 ;
        RECT 22.100 68.400 22.700 79.600 ;
        RECT 22.000 67.600 22.800 68.400 ;
        RECT 23.600 64.200 24.400 75.800 ;
        RECT 25.200 64.200 26.000 77.800 ;
        RECT 26.800 64.200 27.600 77.800 ;
        RECT 33.200 69.600 34.000 70.400 ;
        RECT 44.400 69.600 45.200 70.400 ;
        RECT 49.200 64.200 50.000 77.800 ;
        RECT 50.800 64.200 51.600 77.800 ;
        RECT 52.400 64.200 53.200 75.800 ;
        RECT 54.100 70.400 54.700 81.700 ;
        RECT 54.000 69.600 54.800 70.400 ;
        RECT 54.000 67.600 54.800 68.400 ;
        RECT 55.600 64.200 56.400 75.800 ;
        RECT 58.800 64.200 59.600 75.800 ;
        RECT 60.400 64.200 61.200 77.800 ;
        RECT 62.000 64.200 62.800 77.800 ;
        RECT 63.600 64.200 64.400 77.800 ;
        RECT 73.200 77.600 74.000 78.400 ;
        RECT 76.500 68.400 77.100 93.600 ;
        RECT 81.200 83.600 82.000 84.400 ;
        RECT 81.300 70.400 81.900 83.600 ;
        RECT 82.900 78.400 83.500 95.600 ;
        RECT 86.000 93.600 86.800 94.400 ;
        RECT 87.600 93.600 88.400 94.400 ;
        RECT 90.800 93.600 91.600 94.400 ;
        RECT 86.100 92.400 86.700 93.600 ;
        RECT 87.700 92.400 88.300 93.600 ;
        RECT 90.900 92.400 91.500 93.600 ;
        RECT 98.900 92.400 99.500 95.600 ;
        RECT 100.400 93.600 101.200 94.400 ;
        RECT 100.500 92.400 101.100 93.600 ;
        RECT 86.000 91.600 86.800 92.400 ;
        RECT 87.600 91.600 88.400 92.400 ;
        RECT 90.800 91.600 91.600 92.400 ;
        RECT 98.800 91.600 99.600 92.400 ;
        RECT 100.400 91.600 101.200 92.400 ;
        RECT 90.800 89.600 91.600 90.400 ;
        RECT 82.800 77.600 83.600 78.400 ;
        RECT 90.900 70.400 91.500 89.600 ;
        RECT 92.400 87.600 93.200 88.400 ;
        RECT 95.600 87.600 96.400 88.400 ;
        RECT 94.000 83.600 94.800 84.400 ;
        RECT 94.100 72.400 94.700 83.600 ;
        RECT 94.000 71.600 94.800 72.400 ;
        RECT 95.600 71.600 96.400 72.400 ;
        RECT 95.700 70.400 96.300 71.600 ;
        RECT 81.200 69.600 82.000 70.400 ;
        RECT 84.400 69.600 85.200 70.400 ;
        RECT 90.800 69.600 91.600 70.400 ;
        RECT 95.600 69.600 96.400 70.400 ;
        RECT 74.800 67.600 75.600 68.400 ;
        RECT 76.400 67.600 77.200 68.400 ;
        RECT 86.000 67.600 86.800 68.400 ;
        RECT 86.100 66.400 86.700 67.600 ;
        RECT 81.200 65.600 82.000 66.400 ;
        RECT 86.000 65.600 86.800 66.400 ;
        RECT 81.300 64.400 81.900 65.600 ;
        RECT 81.200 63.600 82.000 64.400 ;
        RECT 87.600 63.600 88.400 64.400 ;
        RECT 4.400 51.600 5.200 52.400 ;
        RECT 4.500 30.400 5.100 51.600 ;
        RECT 9.200 44.200 10.000 57.800 ;
        RECT 10.800 44.200 11.600 57.800 ;
        RECT 12.400 46.200 13.200 57.800 ;
        RECT 14.000 53.600 14.800 54.400 ;
        RECT 15.600 46.200 16.400 57.800 ;
        RECT 18.800 46.200 19.600 57.800 ;
        RECT 20.400 44.200 21.200 57.800 ;
        RECT 22.000 44.200 22.800 57.800 ;
        RECT 23.600 44.200 24.400 57.800 ;
        RECT 57.200 57.600 58.000 58.400 ;
        RECT 68.400 57.600 69.200 58.400 ;
        RECT 42.800 55.000 43.600 55.800 ;
        RECT 44.200 55.000 48.400 55.600 ;
        RECT 49.400 55.000 50.200 55.800 ;
        RECT 52.400 55.600 53.200 56.400 ;
        RECT 34.800 53.600 35.600 54.400 ;
        RECT 41.200 53.600 42.000 54.400 ;
        RECT 42.800 54.200 43.400 55.000 ;
        RECT 44.200 54.800 45.000 55.000 ;
        RECT 47.600 54.800 48.400 55.000 ;
        RECT 42.800 53.600 47.600 54.200 ;
        RECT 34.900 52.400 35.500 53.600 ;
        RECT 34.800 51.600 35.600 52.400 ;
        RECT 41.200 49.600 42.000 50.400 ;
        RECT 42.800 50.200 43.400 53.600 ;
        RECT 46.800 53.400 47.600 53.600 ;
        RECT 49.600 50.200 50.200 55.000 ;
        RECT 50.800 53.600 51.600 54.400 ;
        RECT 50.900 52.400 51.500 53.600 ;
        RECT 50.800 51.600 51.600 52.400 ;
        RECT 52.500 50.400 53.100 55.600 ;
        RECT 55.600 53.600 56.400 54.400 ;
        RECT 57.300 52.400 57.900 57.600 ;
        RECT 68.500 56.400 69.100 57.600 ;
        RECT 65.200 55.600 66.000 56.400 ;
        RECT 68.400 55.600 69.200 56.400 ;
        RECT 73.200 55.600 74.000 56.400 ;
        RECT 81.200 55.600 82.000 56.400 ;
        RECT 84.400 55.600 85.200 56.400 ;
        RECT 81.300 54.400 81.900 55.600 ;
        RECT 66.800 53.600 67.600 54.400 ;
        RECT 71.600 53.600 72.400 54.400 ;
        RECT 76.400 53.600 77.200 54.400 ;
        RECT 81.200 53.600 82.000 54.400 ;
        RECT 71.700 52.400 72.300 53.600 ;
        RECT 57.200 51.600 58.000 52.400 ;
        RECT 58.800 51.600 59.600 52.400 ;
        RECT 71.600 51.600 72.400 52.400 ;
        RECT 81.200 51.600 82.000 52.400 ;
        RECT 81.300 50.400 81.900 51.600 ;
        RECT 4.400 29.600 5.200 30.400 ;
        RECT 9.200 29.600 10.000 30.400 ;
        RECT 4.500 28.400 5.100 29.600 ;
        RECT 4.400 27.600 5.200 28.400 ;
        RECT 4.500 12.400 5.100 27.600 ;
        RECT 14.000 24.200 14.800 37.800 ;
        RECT 15.600 24.200 16.400 37.800 ;
        RECT 17.200 24.200 18.000 35.800 ;
        RECT 18.800 27.600 19.600 28.400 ;
        RECT 20.400 24.200 21.200 35.800 ;
        RECT 23.600 24.200 24.400 35.800 ;
        RECT 25.200 24.200 26.000 37.800 ;
        RECT 26.800 24.200 27.600 37.800 ;
        RECT 28.400 24.200 29.200 37.800 ;
        RECT 41.300 34.400 41.900 49.600 ;
        RECT 42.800 49.400 43.600 50.200 ;
        RECT 49.400 49.400 50.200 50.200 ;
        RECT 52.400 49.600 53.200 50.400 ;
        RECT 63.600 49.600 64.400 50.400 ;
        RECT 81.200 49.600 82.000 50.400 ;
        RECT 84.500 46.400 85.100 55.600 ;
        RECT 87.700 50.400 88.300 63.600 ;
        RECT 89.200 53.600 90.000 54.400 ;
        RECT 89.300 52.400 89.900 53.600 ;
        RECT 89.200 51.600 90.000 52.400 ;
        RECT 90.900 50.400 91.500 69.600 ;
        RECT 94.000 67.600 94.800 68.400 ;
        RECT 94.000 65.600 94.800 66.400 ;
        RECT 94.000 63.600 94.800 64.400 ;
        RECT 94.100 58.400 94.700 63.600 ;
        RECT 94.000 57.600 94.800 58.400 ;
        RECT 100.500 56.300 101.100 91.600 ;
        RECT 102.100 90.400 102.700 95.600 ;
        RECT 105.200 93.600 106.000 94.400 ;
        RECT 105.300 92.400 105.900 93.600 ;
        RECT 106.900 92.400 107.500 95.600 ;
        RECT 105.200 91.600 106.000 92.400 ;
        RECT 106.800 91.600 107.600 92.400 ;
        RECT 102.000 89.600 102.800 90.400 ;
        RECT 103.600 83.600 104.400 84.400 ;
        RECT 103.700 72.400 104.300 83.600 ;
        RECT 103.600 71.600 104.400 72.400 ;
        RECT 103.600 69.600 104.400 70.400 ;
        RECT 100.500 55.700 102.700 56.300 ;
        RECT 102.100 52.400 102.700 55.700 ;
        RECT 92.400 51.600 93.200 52.400 ;
        RECT 97.200 51.600 98.000 52.400 ;
        RECT 102.000 51.600 102.800 52.400 ;
        RECT 87.600 49.600 88.400 50.400 ;
        RECT 90.800 49.600 91.600 50.400 ;
        RECT 87.700 48.400 88.300 49.600 ;
        RECT 87.600 47.600 88.400 48.400 ;
        RECT 90.900 46.400 91.500 49.600 ;
        RECT 92.500 48.400 93.100 51.600 ;
        RECT 92.400 47.600 93.200 48.400 ;
        RECT 84.400 45.600 85.200 46.400 ;
        RECT 90.800 45.600 91.600 46.400 ;
        RECT 52.400 43.600 53.200 44.400 ;
        RECT 58.800 43.600 59.600 44.400 ;
        RECT 70.000 43.600 70.800 44.400 ;
        RECT 49.200 39.600 50.000 40.400 ;
        RECT 41.200 33.600 42.000 34.400 ;
        RECT 30.000 31.600 30.800 32.400 ;
        RECT 30.100 30.400 30.700 31.600 ;
        RECT 30.000 29.600 30.800 30.400 ;
        RECT 46.000 29.600 46.800 30.400 ;
        RECT 39.600 27.600 40.400 28.400 ;
        RECT 49.300 26.400 49.900 39.600 ;
        RECT 52.500 30.400 53.100 43.600 ;
        RECT 58.900 42.400 59.500 43.600 ;
        RECT 58.800 41.600 59.600 42.400 ;
        RECT 58.900 40.400 59.500 41.600 ;
        RECT 70.100 40.400 70.700 43.600 ;
        RECT 58.800 39.600 59.600 40.400 ;
        RECT 63.600 39.600 64.400 40.400 ;
        RECT 70.000 39.600 70.800 40.400 ;
        RECT 54.000 31.600 54.800 32.400 ;
        RECT 54.100 30.400 54.700 31.600 ;
        RECT 52.400 29.600 53.200 30.400 ;
        RECT 54.000 29.600 54.800 30.400 ;
        RECT 55.600 29.600 56.400 30.400 ;
        RECT 50.800 27.600 51.600 28.400 ;
        RECT 49.200 25.600 50.000 26.400 ;
        RECT 4.400 11.600 5.200 12.400 ;
        RECT 9.200 4.200 10.000 17.800 ;
        RECT 10.800 4.200 11.600 17.800 ;
        RECT 12.400 6.200 13.200 17.800 ;
        RECT 14.000 13.600 14.800 14.400 ;
        RECT 15.600 6.200 16.400 17.800 ;
        RECT 18.800 6.200 19.600 17.800 ;
        RECT 20.400 4.200 21.200 17.800 ;
        RECT 22.000 4.200 22.800 17.800 ;
        RECT 23.600 4.200 24.400 17.800 ;
        RECT 41.200 15.600 42.000 16.400 ;
        RECT 41.300 14.400 41.900 15.600 ;
        RECT 42.800 15.000 43.600 15.800 ;
        RECT 44.200 15.000 48.400 15.600 ;
        RECT 49.400 15.000 50.200 15.800 ;
        RECT 34.800 13.600 35.600 14.400 ;
        RECT 41.200 13.600 42.000 14.400 ;
        RECT 42.800 14.200 43.400 15.000 ;
        RECT 44.200 14.800 45.000 15.000 ;
        RECT 47.600 14.800 48.400 15.000 ;
        RECT 42.800 13.600 47.600 14.200 ;
        RECT 34.900 12.400 35.500 13.600 ;
        RECT 34.800 11.600 35.600 12.400 ;
        RECT 42.800 10.200 43.400 13.600 ;
        RECT 46.800 13.400 47.600 13.600 ;
        RECT 49.600 10.200 50.200 15.000 ;
        RECT 50.900 14.400 51.500 27.600 ;
        RECT 50.800 13.600 51.600 14.400 ;
        RECT 55.700 12.400 56.300 29.600 ;
        RECT 58.800 24.200 59.600 37.800 ;
        RECT 60.400 24.200 61.200 37.800 ;
        RECT 62.000 24.200 62.800 35.800 ;
        RECT 63.700 28.400 64.300 39.600 ;
        RECT 63.600 27.600 64.400 28.400 ;
        RECT 65.200 24.200 66.000 35.800 ;
        RECT 68.400 24.200 69.200 35.800 ;
        RECT 70.000 24.200 70.800 37.800 ;
        RECT 71.600 24.200 72.400 37.800 ;
        RECT 73.200 24.200 74.000 37.800 ;
        RECT 84.500 34.400 85.100 45.600 ;
        RECT 89.200 43.600 90.000 44.400 ;
        RECT 84.400 33.600 85.200 34.400 ;
        RECT 89.300 32.400 89.900 43.600 ;
        RECT 92.400 41.600 93.200 42.400 ;
        RECT 92.500 34.400 93.100 41.600 ;
        RECT 92.400 33.600 93.200 34.400 ;
        RECT 89.200 31.600 90.000 32.400 ;
        RECT 95.600 31.600 96.400 32.400 ;
        RECT 103.600 31.600 104.400 32.400 ;
        RECT 89.300 28.400 89.900 31.600 ;
        RECT 94.000 29.600 94.800 30.400 ;
        RECT 89.200 27.600 90.000 28.400 ;
        RECT 94.000 27.600 94.800 28.400 ;
        RECT 86.000 25.600 86.800 26.400 ;
        RECT 89.200 25.600 90.000 26.400 ;
        RECT 55.600 11.600 56.400 12.400 ;
        RECT 42.800 9.400 43.600 10.200 ;
        RECT 49.400 9.400 50.200 10.200 ;
        RECT 60.400 4.200 61.200 17.800 ;
        RECT 62.000 4.200 62.800 17.800 ;
        RECT 63.600 6.200 64.400 17.800 ;
        RECT 65.200 13.600 66.000 14.400 ;
        RECT 66.800 6.200 67.600 17.800 ;
        RECT 70.000 6.200 70.800 17.800 ;
        RECT 71.600 4.200 72.400 17.800 ;
        RECT 73.200 4.200 74.000 17.800 ;
        RECT 74.800 4.200 75.600 17.800 ;
        RECT 86.100 16.400 86.700 25.600 ;
        RECT 89.300 16.400 89.900 25.600 ;
        RECT 92.400 23.600 93.200 24.400 ;
        RECT 86.000 15.600 86.800 16.400 ;
        RECT 89.200 15.600 90.000 16.400 ;
        RECT 92.500 10.400 93.100 23.600 ;
        RECT 94.100 18.400 94.700 27.600 ;
        RECT 94.000 17.600 94.800 18.400 ;
        RECT 95.700 16.400 96.300 31.600 ;
        RECT 97.200 29.600 98.000 30.400 ;
        RECT 100.400 29.600 101.200 30.400 ;
        RECT 98.800 25.600 99.600 26.400 ;
        RECT 100.500 16.400 101.100 29.600 ;
        RECT 95.600 15.600 96.400 16.400 ;
        RECT 100.400 15.600 101.200 16.400 ;
        RECT 95.600 13.600 96.400 14.400 ;
        RECT 98.800 13.600 99.600 14.400 ;
        RECT 103.700 12.400 104.300 31.600 ;
        RECT 105.200 29.600 106.000 30.400 ;
        RECT 105.300 26.400 105.900 29.600 ;
        RECT 105.200 25.600 106.000 26.400 ;
        RECT 108.400 25.600 109.200 26.400 ;
        RECT 106.800 13.600 107.600 14.400 ;
        RECT 103.600 11.600 104.400 12.400 ;
        RECT 108.500 10.400 109.100 25.600 ;
        RECT 92.400 9.600 93.200 10.400 ;
        RECT 95.600 9.600 96.400 10.400 ;
        RECT 108.400 9.600 109.200 10.400 ;
      LAYER metal3 ;
        RECT 20.400 96.300 21.200 96.400 ;
        RECT 76.400 96.300 77.200 96.400 ;
        RECT 20.400 95.700 77.200 96.300 ;
        RECT 20.400 95.600 21.200 95.700 ;
        RECT 76.400 95.600 77.200 95.700 ;
        RECT 82.800 96.300 83.600 96.400 ;
        RECT 98.800 96.300 99.600 96.400 ;
        RECT 102.000 96.300 102.800 96.400 ;
        RECT 106.800 96.300 107.600 96.400 ;
        RECT 82.800 95.700 107.600 96.300 ;
        RECT 82.800 95.600 83.600 95.700 ;
        RECT 98.800 95.600 99.600 95.700 ;
        RECT 102.000 95.600 102.800 95.700 ;
        RECT 106.800 95.600 107.600 95.700 ;
        RECT 6.000 94.300 6.800 94.400 ;
        RECT 15.600 94.300 16.400 94.400 ;
        RECT 87.600 94.300 88.400 94.400 ;
        RECT 90.800 94.300 91.600 94.400 ;
        RECT 6.000 93.700 91.600 94.300 ;
        RECT 6.000 93.600 6.800 93.700 ;
        RECT 15.600 93.600 16.400 93.700 ;
        RECT 87.600 93.600 88.400 93.700 ;
        RECT 90.800 93.600 91.600 93.700 ;
        RECT 2.800 92.300 3.600 92.400 ;
        RECT 7.600 92.300 8.400 92.400 ;
        RECT 22.000 92.300 22.800 92.400 ;
        RECT 2.800 91.700 22.800 92.300 ;
        RECT 2.800 91.600 3.600 91.700 ;
        RECT 7.600 91.600 8.400 91.700 ;
        RECT 22.000 91.600 22.800 91.700 ;
        RECT 44.400 92.300 45.200 92.400 ;
        RECT 65.200 92.300 66.000 92.400 ;
        RECT 44.400 91.700 66.000 92.300 ;
        RECT 44.400 91.600 45.200 91.700 ;
        RECT 65.200 91.600 66.000 91.700 ;
        RECT 66.800 92.300 67.600 92.400 ;
        RECT 86.000 92.300 86.800 92.400 ;
        RECT 100.400 92.300 101.200 92.400 ;
        RECT 105.200 92.300 106.000 92.400 ;
        RECT 66.800 91.700 106.000 92.300 ;
        RECT 66.800 91.600 67.600 91.700 ;
        RECT 86.000 91.600 86.800 91.700 ;
        RECT 100.400 91.600 101.200 91.700 ;
        RECT 105.200 91.600 106.000 91.700 ;
        RECT 92.400 88.300 93.200 88.400 ;
        RECT 95.600 88.300 96.400 88.400 ;
        RECT 92.400 87.700 96.400 88.300 ;
        RECT 92.400 87.600 93.200 87.700 ;
        RECT 95.600 87.600 96.400 87.700 ;
        RECT 15.600 80.300 16.400 80.400 ;
        RECT 22.000 80.300 22.800 80.400 ;
        RECT 15.600 79.700 22.800 80.300 ;
        RECT 15.600 79.600 16.400 79.700 ;
        RECT 22.000 79.600 22.800 79.700 ;
        RECT 73.200 78.300 74.000 78.400 ;
        RECT 82.800 78.300 83.600 78.400 ;
        RECT 73.200 77.700 83.600 78.300 ;
        RECT 73.200 77.600 74.000 77.700 ;
        RECT 82.800 77.600 83.600 77.700 ;
        RECT 58.800 72.300 59.600 72.400 ;
        RECT 94.000 72.300 94.800 72.400 ;
        RECT 58.800 71.700 94.800 72.300 ;
        RECT 58.800 71.600 59.600 71.700 ;
        RECT 94.000 71.600 94.800 71.700 ;
        RECT 95.600 72.300 96.400 72.400 ;
        RECT 103.600 72.300 104.400 72.400 ;
        RECT 95.600 71.700 104.400 72.300 ;
        RECT 95.600 71.600 96.400 71.700 ;
        RECT 103.600 71.600 104.400 71.700 ;
        RECT 4.400 70.300 5.200 70.400 ;
        RECT 10.800 70.300 11.600 70.400 ;
        RECT 4.400 69.700 11.600 70.300 ;
        RECT 4.400 69.600 5.200 69.700 ;
        RECT 10.800 69.600 11.600 69.700 ;
        RECT 33.200 70.300 34.000 70.400 ;
        RECT 44.400 70.300 45.200 70.400 ;
        RECT 33.200 69.700 45.200 70.300 ;
        RECT 33.200 69.600 34.000 69.700 ;
        RECT 44.400 69.600 45.200 69.700 ;
        RECT 81.200 70.300 82.000 70.400 ;
        RECT 84.400 70.300 85.200 70.400 ;
        RECT 81.200 69.700 85.200 70.300 ;
        RECT 81.200 69.600 82.000 69.700 ;
        RECT 84.400 69.600 85.200 69.700 ;
        RECT 90.800 70.300 91.600 70.400 ;
        RECT 103.600 70.300 104.400 70.400 ;
        RECT 90.800 69.700 104.400 70.300 ;
        RECT 90.800 69.600 91.600 69.700 ;
        RECT 103.600 69.600 104.400 69.700 ;
        RECT 54.000 68.300 54.800 68.400 ;
        RECT 74.800 68.300 75.600 68.400 ;
        RECT 54.000 67.700 75.600 68.300 ;
        RECT 54.000 67.600 54.800 67.700 ;
        RECT 74.800 67.600 75.600 67.700 ;
        RECT 76.400 68.300 77.200 68.400 ;
        RECT 86.000 68.300 86.800 68.400 ;
        RECT 94.000 68.300 94.800 68.400 ;
        RECT 76.400 67.700 94.800 68.300 ;
        RECT 76.400 67.600 77.200 67.700 ;
        RECT 86.000 67.600 86.800 67.700 ;
        RECT 94.000 67.600 94.800 67.700 ;
        RECT 94.000 65.600 94.800 66.400 ;
        RECT 81.200 64.300 82.000 64.400 ;
        RECT 87.600 64.300 88.400 64.400 ;
        RECT 81.200 63.700 88.400 64.300 ;
        RECT 81.200 63.600 82.000 63.700 ;
        RECT 87.600 63.600 88.400 63.700 ;
        RECT 57.200 58.300 58.000 58.400 ;
        RECT 68.400 58.300 69.200 58.400 ;
        RECT 94.000 58.300 94.800 58.400 ;
        RECT 57.200 57.700 94.800 58.300 ;
        RECT 57.200 57.600 58.000 57.700 ;
        RECT 68.400 57.600 69.200 57.700 ;
        RECT 94.000 57.600 94.800 57.700 ;
        RECT 65.200 56.300 66.000 56.400 ;
        RECT 73.200 56.300 74.000 56.400 ;
        RECT 65.200 55.700 74.000 56.300 ;
        RECT 65.200 55.600 66.000 55.700 ;
        RECT 73.200 55.600 74.000 55.700 ;
        RECT 14.000 54.300 14.800 54.400 ;
        RECT 34.800 54.300 35.600 54.400 ;
        RECT 14.000 53.700 35.600 54.300 ;
        RECT 14.000 53.600 14.800 53.700 ;
        RECT 34.800 53.600 35.600 53.700 ;
        RECT 41.200 54.300 42.000 54.400 ;
        RECT 55.600 54.300 56.400 54.400 ;
        RECT 66.800 54.300 67.600 54.400 ;
        RECT 41.200 53.700 67.600 54.300 ;
        RECT 41.200 53.600 42.000 53.700 ;
        RECT 55.600 53.600 56.400 53.700 ;
        RECT 66.800 53.600 67.600 53.700 ;
        RECT 71.600 54.300 72.400 54.400 ;
        RECT 76.400 54.300 77.200 54.400 ;
        RECT 71.600 53.700 77.200 54.300 ;
        RECT 71.600 53.600 72.400 53.700 ;
        RECT 76.400 53.600 77.200 53.700 ;
        RECT 81.200 54.300 82.000 54.400 ;
        RECT 89.200 54.300 90.000 54.400 ;
        RECT 81.200 53.700 90.000 54.300 ;
        RECT 81.200 53.600 82.000 53.700 ;
        RECT 89.200 53.600 90.000 53.700 ;
        RECT 50.800 52.300 51.600 52.400 ;
        RECT 58.800 52.300 59.600 52.400 ;
        RECT 50.800 51.700 59.600 52.300 ;
        RECT 66.900 52.300 67.500 53.600 ;
        RECT 97.200 52.300 98.000 52.400 ;
        RECT 66.900 51.700 98.000 52.300 ;
        RECT 50.800 51.600 51.600 51.700 ;
        RECT 58.800 51.600 59.600 51.700 ;
        RECT 97.200 51.600 98.000 51.700 ;
        RECT 41.200 50.300 42.000 50.400 ;
        RECT 52.400 50.300 53.200 50.400 ;
        RECT 63.600 50.300 64.400 50.400 ;
        RECT 41.200 49.700 64.400 50.300 ;
        RECT 41.200 49.600 42.000 49.700 ;
        RECT 52.400 49.600 53.200 49.700 ;
        RECT 63.600 49.600 64.400 49.700 ;
        RECT 81.200 50.300 82.000 50.400 ;
        RECT 87.600 50.300 88.400 50.400 ;
        RECT 81.200 49.700 88.400 50.300 ;
        RECT 81.200 49.600 82.000 49.700 ;
        RECT 87.600 49.600 88.400 49.700 ;
        RECT 63.700 48.300 64.300 49.600 ;
        RECT 92.400 48.300 93.200 48.400 ;
        RECT 63.700 47.700 93.200 48.300 ;
        RECT 92.400 47.600 93.200 47.700 ;
        RECT 84.400 46.300 85.200 46.400 ;
        RECT 90.800 46.300 91.600 46.400 ;
        RECT 84.400 45.700 91.600 46.300 ;
        RECT 84.400 45.600 85.200 45.700 ;
        RECT 90.800 45.600 91.600 45.700 ;
        RECT 58.800 42.300 59.600 42.400 ;
        RECT 92.400 42.300 93.200 42.400 ;
        RECT 58.800 41.700 93.200 42.300 ;
        RECT 58.800 41.600 59.600 41.700 ;
        RECT 92.400 41.600 93.200 41.700 ;
        RECT 49.200 40.300 50.000 40.400 ;
        RECT 58.800 40.300 59.600 40.400 ;
        RECT 49.200 39.700 59.600 40.300 ;
        RECT 49.200 39.600 50.000 39.700 ;
        RECT 58.800 39.600 59.600 39.700 ;
        RECT 63.600 40.300 64.400 40.400 ;
        RECT 70.000 40.300 70.800 40.400 ;
        RECT 63.600 39.700 70.800 40.300 ;
        RECT 63.600 39.600 64.400 39.700 ;
        RECT 70.000 39.600 70.800 39.700 ;
        RECT 30.000 32.300 30.800 32.400 ;
        RECT 54.000 32.300 54.800 32.400 ;
        RECT 30.000 31.700 54.800 32.300 ;
        RECT 30.000 31.600 30.800 31.700 ;
        RECT 54.000 31.600 54.800 31.700 ;
        RECT 89.200 32.300 90.000 32.400 ;
        RECT 103.600 32.300 104.400 32.400 ;
        RECT 89.200 31.700 104.400 32.300 ;
        RECT 89.200 31.600 90.000 31.700 ;
        RECT 103.600 31.600 104.400 31.700 ;
        RECT 4.400 30.300 5.200 30.400 ;
        RECT 9.200 30.300 10.000 30.400 ;
        RECT 4.400 29.700 10.000 30.300 ;
        RECT 4.400 29.600 5.200 29.700 ;
        RECT 9.200 29.600 10.000 29.700 ;
        RECT 46.000 30.300 46.800 30.400 ;
        RECT 52.400 30.300 53.200 30.400 ;
        RECT 46.000 29.700 53.200 30.300 ;
        RECT 46.000 29.600 46.800 29.700 ;
        RECT 52.400 29.600 53.200 29.700 ;
        RECT 94.000 30.300 94.800 30.400 ;
        RECT 97.200 30.300 98.000 30.400 ;
        RECT 94.000 29.700 98.000 30.300 ;
        RECT 94.000 29.600 94.800 29.700 ;
        RECT 97.200 29.600 98.000 29.700 ;
        RECT 18.800 28.300 19.600 28.400 ;
        RECT 39.600 28.300 40.400 28.400 ;
        RECT 18.800 27.700 40.400 28.300 ;
        RECT 18.800 27.600 19.600 27.700 ;
        RECT 39.600 27.600 40.400 27.700 ;
        RECT 50.800 28.300 51.600 28.400 ;
        RECT 89.200 28.300 90.000 28.400 ;
        RECT 50.800 27.700 90.000 28.300 ;
        RECT 50.800 27.600 51.600 27.700 ;
        RECT 89.200 27.600 90.000 27.700 ;
        RECT 94.000 27.600 94.800 28.400 ;
        RECT 86.000 26.300 86.800 26.400 ;
        RECT 98.800 26.300 99.600 26.400 ;
        RECT 105.200 26.300 106.000 26.400 ;
        RECT 108.400 26.300 109.200 26.400 ;
        RECT 86.000 25.700 109.200 26.300 ;
        RECT 86.000 25.600 86.800 25.700 ;
        RECT 98.800 25.600 99.600 25.700 ;
        RECT 105.200 25.600 106.000 25.700 ;
        RECT 108.400 25.600 109.200 25.700 ;
        RECT 41.200 16.300 42.000 16.400 ;
        RECT 95.600 16.300 96.400 16.400 ;
        RECT 100.400 16.300 101.200 16.400 ;
        RECT 41.200 15.700 101.200 16.300 ;
        RECT 41.200 15.600 42.000 15.700 ;
        RECT 95.600 15.600 96.400 15.700 ;
        RECT 100.400 15.600 101.200 15.700 ;
        RECT 14.000 14.300 14.800 14.400 ;
        RECT 34.800 14.300 35.600 14.400 ;
        RECT 14.000 13.700 35.600 14.300 ;
        RECT 14.000 13.600 14.800 13.700 ;
        RECT 34.800 13.600 35.600 13.700 ;
        RECT 65.200 14.300 66.000 14.400 ;
        RECT 95.600 14.300 96.400 14.400 ;
        RECT 65.200 13.700 96.400 14.300 ;
        RECT 65.200 13.600 66.000 13.700 ;
        RECT 95.600 13.600 96.400 13.700 ;
        RECT 98.800 14.300 99.600 14.400 ;
        RECT 106.800 14.300 107.600 14.400 ;
        RECT 98.800 13.700 107.600 14.300 ;
        RECT 98.800 13.600 99.600 13.700 ;
        RECT 106.800 13.600 107.600 13.700 ;
        RECT 92.400 10.300 93.200 10.400 ;
        RECT 95.600 10.300 96.400 10.400 ;
        RECT 92.400 9.700 96.400 10.300 ;
        RECT 92.400 9.600 93.200 9.700 ;
        RECT 95.600 9.600 96.400 9.700 ;
      LAYER metal4 ;
        RECT 58.600 51.400 59.800 72.600 ;
        RECT 93.800 27.400 95.000 66.600 ;
  END
END up_counter
END LIBRARY

