magic
tech scmos
magscale 1 2
timestamp 1733888598
<< metal1 >>
rect 792 1006 798 1014
rect 806 1006 812 1014
rect 820 1006 826 1014
rect 834 1006 840 1014
rect 253 977 300 983
rect 125 943 131 963
rect 196 956 204 964
rect 93 937 131 943
rect 638 937 668 943
rect 12 924 20 928
rect 205 917 220 923
rect 205 897 211 917
rect 660 917 712 923
rect 893 897 908 903
rect 820 837 835 843
rect 344 806 350 814
rect 358 806 364 814
rect 372 806 378 814
rect 386 806 392 814
rect 893 697 956 703
rect 756 677 835 683
rect 1069 677 1100 683
rect 792 606 798 614
rect 806 606 812 614
rect 820 606 826 614
rect 834 606 840 614
rect 1053 577 1084 583
rect 621 557 652 563
rect 749 557 812 563
rect 334 537 412 543
rect 772 537 835 543
rect 356 517 451 523
rect 708 436 710 444
rect 344 406 350 414
rect 358 406 364 414
rect 372 406 378 414
rect 386 406 392 414
rect 381 337 412 343
rect 829 337 844 343
rect 29 277 44 283
rect 404 277 483 283
rect 1085 277 1100 283
rect 829 257 892 263
rect 792 206 798 214
rect 806 206 812 214
rect 820 206 826 214
rect 834 206 840 214
rect 845 157 860 163
rect 900 157 931 163
rect 334 137 412 143
rect 964 137 979 143
rect 1021 137 1043 143
rect 356 117 451 123
rect 1044 117 1059 123
rect 344 6 350 14
rect 358 6 364 14
rect 372 6 378 14
rect 386 6 392 14
<< m2contact >>
rect 798 1006 806 1014
rect 812 1006 820 1014
rect 826 1006 834 1014
rect 300 976 308 984
rect 108 956 116 964
rect 204 956 212 964
rect 476 956 484 964
rect 828 956 836 964
rect 172 936 180 944
rect 444 936 452 944
rect 668 936 676 944
rect 764 936 772 944
rect 860 936 868 944
rect 1004 936 1012 944
rect 1052 936 1060 944
rect 12 916 20 924
rect 28 916 36 924
rect 60 916 68 924
rect 76 916 84 924
rect 156 916 164 924
rect 220 916 228 924
rect 556 916 564 924
rect 652 916 660 924
rect 876 916 884 924
rect 908 916 916 924
rect 988 916 996 924
rect 1068 916 1076 924
rect 380 900 388 908
rect 908 896 916 904
rect 1020 896 1028 904
rect 924 876 932 884
rect 956 876 964 884
rect 1100 876 1108 884
rect 380 854 388 862
rect 156 836 164 844
rect 812 836 820 844
rect 940 836 948 844
rect 1036 836 1044 844
rect 350 806 358 814
rect 364 806 372 814
rect 378 806 386 814
rect 28 776 36 784
rect 316 776 324 784
rect 444 776 452 784
rect 732 776 740 784
rect 316 716 324 724
rect 444 716 452 724
rect 108 696 116 704
rect 332 696 340 704
rect 444 696 452 704
rect 540 696 548 704
rect 844 696 852 704
rect 956 696 964 704
rect 1036 696 1044 704
rect 220 676 228 684
rect 540 676 548 684
rect 748 676 756 684
rect 940 676 948 684
rect 1100 676 1108 684
rect 188 656 196 664
rect 572 656 580 664
rect 812 656 820 664
rect 860 656 868 664
rect 940 656 948 664
rect 876 636 884 644
rect 940 636 948 644
rect 798 606 806 614
rect 812 606 820 614
rect 826 606 834 614
rect 1084 576 1092 584
rect 172 556 180 564
rect 524 556 532 564
rect 652 556 660 564
rect 684 556 692 564
rect 732 556 740 564
rect 812 556 820 564
rect 844 556 852 564
rect 140 536 148 544
rect 412 536 420 544
rect 508 536 516 544
rect 556 536 564 544
rect 668 536 676 544
rect 764 536 772 544
rect 1004 536 1012 544
rect 44 516 52 524
rect 348 516 356 524
rect 572 516 580 524
rect 588 516 596 524
rect 716 516 724 524
rect 812 516 820 524
rect 892 516 900 524
rect 924 516 932 524
rect 972 516 980 524
rect 1020 516 1028 524
rect 76 500 84 508
rect 636 496 644 504
rect 908 496 916 504
rect 876 476 884 484
rect 956 476 964 484
rect 76 436 84 444
rect 524 436 532 444
rect 588 436 596 444
rect 700 436 708 444
rect 892 436 900 444
rect 350 406 358 414
rect 364 406 372 414
rect 378 406 386 414
rect 92 376 100 384
rect 572 358 580 366
rect 412 336 420 344
rect 844 336 852 344
rect 924 336 932 344
rect 1036 336 1044 344
rect 92 316 100 324
rect 572 312 580 320
rect 956 316 964 324
rect 92 296 100 304
rect 300 296 308 304
rect 460 296 468 304
rect 540 296 548 304
rect 556 296 564 304
rect 940 296 948 304
rect 972 296 980 304
rect 1004 296 1012 304
rect 1052 296 1060 304
rect 12 276 20 284
rect 44 276 52 284
rect 188 276 196 284
rect 396 276 404 284
rect 636 276 644 284
rect 1100 276 1108 284
rect 220 256 228 264
rect 492 256 500 264
rect 668 256 676 264
rect 892 256 900 264
rect 988 256 996 264
rect 924 236 932 244
rect 798 206 806 214
rect 812 206 820 214
rect 826 206 834 214
rect 940 176 948 184
rect 172 156 180 164
rect 684 156 692 164
rect 860 156 868 164
rect 892 156 900 164
rect 1004 156 1012 164
rect 140 136 148 144
rect 412 136 420 144
rect 508 136 516 144
rect 652 136 660 144
rect 956 136 964 144
rect 988 136 996 144
rect 1068 136 1076 144
rect 44 116 52 124
rect 348 116 356 124
rect 556 116 564 124
rect 1036 116 1044 124
rect 44 96 52 104
rect 556 96 564 104
rect 956 96 964 104
rect 1084 96 1092 104
rect 44 36 52 44
rect 556 36 564 44
rect 350 6 358 14
rect 364 6 372 14
rect 378 6 386 14
<< metal2 >>
rect 792 1006 798 1014
rect 806 1006 812 1014
rect 820 1006 826 1014
rect 834 1006 840 1014
rect 61 924 67 936
rect 13 904 19 916
rect 29 784 35 916
rect 109 904 115 956
rect 157 924 163 936
rect 173 904 179 936
rect 445 924 451 936
rect 381 862 387 900
rect 157 804 163 836
rect 344 806 350 814
rect 358 806 364 814
rect 372 806 378 814
rect 386 806 392 814
rect 45 524 51 696
rect 221 684 227 796
rect 317 724 323 776
rect 445 724 451 776
rect 477 664 483 956
rect 765 944 771 956
rect 669 924 675 936
rect 557 823 563 916
rect 541 817 563 823
rect 541 704 547 817
rect 765 684 771 936
rect 813 704 819 836
rect 829 784 835 956
rect 861 924 867 936
rect 877 924 883 936
rect 909 924 915 936
rect 989 924 995 956
rect 1005 924 1011 936
rect 909 704 915 896
rect 941 724 947 836
rect 957 704 963 716
rect 861 664 867 676
rect 189 603 195 656
rect 813 644 819 656
rect 792 606 798 614
rect 806 606 812 614
rect 820 606 826 614
rect 834 606 840 614
rect 173 597 195 603
rect 173 564 179 597
rect 45 304 51 516
rect 77 444 83 500
rect 173 384 179 556
rect 349 524 355 536
rect 509 524 515 536
rect 525 504 531 556
rect 573 524 579 576
rect 685 564 691 576
rect 813 544 819 556
rect 717 524 723 536
rect 813 504 819 516
rect 344 406 350 414
rect 358 406 364 414
rect 372 406 378 414
rect 386 406 392 414
rect 93 324 99 376
rect 221 324 227 376
rect 413 344 419 496
rect 845 464 851 556
rect 877 504 883 636
rect 893 524 899 536
rect 909 504 915 696
rect 941 584 947 636
rect 1005 563 1011 916
rect 1021 904 1027 956
rect 1053 924 1059 936
rect 1069 924 1075 956
rect 1037 724 1043 836
rect 1085 584 1091 936
rect 1101 884 1107 896
rect 1101 684 1107 696
rect 1005 557 1027 563
rect 1021 524 1027 557
rect 877 484 883 496
rect 909 464 915 496
rect 925 484 931 516
rect 957 484 963 496
rect 45 284 51 296
rect 45 124 51 276
rect 221 264 227 316
rect 301 304 307 316
rect 493 264 499 396
rect 525 304 531 436
rect 589 424 595 436
rect 589 404 595 416
rect 701 404 707 436
rect 573 320 579 358
rect 541 304 547 316
rect 221 204 227 256
rect 173 164 179 196
rect 413 144 419 156
rect 509 144 515 276
rect 349 124 355 136
rect 557 124 563 296
rect 637 284 643 396
rect 845 344 851 456
rect 893 324 899 436
rect 925 344 931 416
rect 893 284 899 316
rect 669 204 675 256
rect 792 206 798 214
rect 806 206 812 214
rect 820 206 826 214
rect 834 206 840 214
rect 685 164 691 196
rect 861 164 867 256
rect 893 164 899 256
rect 925 104 931 236
rect 941 184 947 276
rect 957 164 963 316
rect 1005 164 1011 296
rect 1037 124 1043 316
rect 1053 264 1059 296
rect 1101 284 1107 296
rect 1085 104 1091 256
rect 45 44 51 96
rect 557 44 563 96
rect 344 6 350 14
rect 358 6 364 14
rect 372 6 378 14
rect 386 6 392 14
<< m3contact >>
rect 798 1006 806 1014
rect 812 1006 820 1014
rect 826 1006 834 1014
rect 300 976 308 984
rect 204 956 212 964
rect 764 956 772 964
rect 828 956 836 964
rect 988 956 996 964
rect 1020 956 1028 964
rect 1068 956 1076 964
rect 60 936 68 944
rect 28 916 36 924
rect 76 916 84 924
rect 12 896 20 904
rect 156 936 164 944
rect 220 916 228 924
rect 444 916 452 924
rect 108 896 116 904
rect 172 896 180 904
rect 350 806 358 814
rect 364 806 372 814
rect 378 806 386 814
rect 156 796 164 804
rect 220 796 228 804
rect 44 696 52 704
rect 108 696 116 704
rect 332 696 340 704
rect 444 696 452 704
rect 652 916 660 924
rect 668 916 676 924
rect 732 776 740 784
rect 876 936 884 944
rect 908 936 916 944
rect 860 916 868 924
rect 1004 916 1012 924
rect 828 776 836 784
rect 924 876 932 884
rect 956 876 964 884
rect 940 716 948 724
rect 956 716 964 724
rect 812 696 820 704
rect 844 696 852 704
rect 908 696 916 704
rect 540 676 548 684
rect 748 676 756 684
rect 764 676 772 684
rect 860 676 868 684
rect 188 656 196 664
rect 476 656 484 664
rect 572 656 580 664
rect 812 636 820 644
rect 876 636 884 644
rect 798 606 806 614
rect 812 606 820 614
rect 826 606 834 614
rect 572 576 580 584
rect 684 576 692 584
rect 140 536 148 544
rect 348 536 356 544
rect 412 536 420 544
rect 508 516 516 524
rect 556 536 564 544
rect 652 556 660 564
rect 732 556 740 564
rect 668 536 676 544
rect 716 536 724 544
rect 764 536 772 544
rect 812 536 820 544
rect 588 516 596 524
rect 412 496 420 504
rect 524 496 532 504
rect 636 496 644 504
rect 812 496 820 504
rect 350 406 358 414
rect 364 406 372 414
rect 378 406 386 414
rect 172 376 180 384
rect 220 376 228 384
rect 892 536 900 544
rect 940 676 948 684
rect 940 656 948 664
rect 940 576 948 584
rect 1084 936 1092 944
rect 1052 916 1060 924
rect 1036 716 1044 724
rect 1036 696 1044 704
rect 1100 896 1108 904
rect 1100 696 1108 704
rect 1004 536 1012 544
rect 972 516 980 524
rect 876 496 884 504
rect 956 496 964 504
rect 924 476 932 484
rect 844 456 852 464
rect 908 456 916 464
rect 492 396 500 404
rect 220 316 228 324
rect 300 316 308 324
rect 44 296 52 304
rect 92 296 100 304
rect 12 276 20 284
rect 188 276 196 284
rect 460 296 468 304
rect 396 276 404 284
rect 588 416 596 424
rect 588 396 596 404
rect 636 396 644 404
rect 700 396 708 404
rect 540 316 548 324
rect 524 296 532 304
rect 508 276 516 284
rect 172 196 180 204
rect 220 196 228 204
rect 412 156 420 164
rect 140 136 148 144
rect 348 136 356 144
rect 924 416 932 424
rect 1036 336 1044 344
rect 892 316 900 324
rect 1036 316 1044 324
rect 940 296 948 304
rect 892 276 900 284
rect 940 276 948 284
rect 860 256 868 264
rect 798 206 806 214
rect 812 206 820 214
rect 826 206 834 214
rect 668 196 676 204
rect 684 196 692 204
rect 652 136 660 144
rect 972 296 980 304
rect 988 256 996 264
rect 956 156 964 164
rect 1004 156 1012 164
rect 956 136 964 144
rect 988 136 996 144
rect 1100 296 1108 304
rect 1052 256 1060 264
rect 1084 256 1092 264
rect 1068 136 1076 144
rect 924 96 932 104
rect 956 96 964 104
rect 350 6 358 14
rect 364 6 372 14
rect 378 6 386 14
<< metal3 >>
rect 792 1014 840 1016
rect 792 1006 796 1014
rect 806 1006 812 1014
rect 820 1006 826 1014
rect 836 1006 840 1014
rect 792 1004 840 1006
rect 308 977 1139 983
rect 212 957 764 963
rect 836 957 988 963
rect 996 957 1020 963
rect 1028 957 1068 963
rect 68 937 156 943
rect 164 937 876 943
rect 884 937 908 943
rect 1092 937 1139 943
rect 36 917 76 923
rect 84 917 220 923
rect 452 917 652 923
rect 676 917 860 923
rect 868 917 1004 923
rect 1012 917 1052 923
rect -19 897 12 903
rect 20 897 108 903
rect 116 897 172 903
rect 1108 897 1139 903
rect 932 877 956 883
rect 344 814 392 816
rect 344 806 348 814
rect 358 806 364 814
rect 372 806 378 814
rect 388 806 392 814
rect 344 804 392 806
rect 164 797 220 803
rect 740 777 828 783
rect 596 717 940 723
rect 964 717 1036 723
rect 52 697 108 703
rect 340 697 444 703
rect 820 697 844 703
rect 916 697 1036 703
rect 1108 697 1139 703
rect 548 677 748 683
rect 772 677 860 683
rect 868 677 940 683
rect 196 657 476 663
rect 484 657 572 663
rect 820 637 876 643
rect 792 614 840 616
rect 792 606 796 614
rect 806 606 812 614
rect 820 606 826 614
rect 836 606 840 614
rect 792 604 840 606
rect 580 577 684 583
rect 692 577 940 583
rect 660 557 732 563
rect 148 537 348 543
rect 420 537 556 543
rect 564 537 668 543
rect 724 537 764 543
rect 820 537 892 543
rect 1012 537 1139 543
rect 516 517 588 523
rect 669 523 675 536
rect 669 517 972 523
rect 420 497 524 503
rect 532 497 636 503
rect 820 497 876 503
rect 964 497 1139 503
rect 637 483 643 496
rect 637 477 924 483
rect 852 457 908 463
rect 596 417 924 423
rect 344 414 392 416
rect 344 406 348 414
rect 358 406 364 414
rect 372 406 378 414
rect 388 406 392 414
rect 344 404 392 406
rect 500 397 588 403
rect 644 397 700 403
rect 180 377 220 383
rect 1044 337 1139 343
rect -19 317 220 323
rect 308 317 540 323
rect 900 317 1036 323
rect 52 297 92 303
rect 468 297 524 303
rect 948 297 972 303
rect 1108 297 1139 303
rect -19 277 12 283
rect 196 277 396 283
rect 516 277 892 283
rect 868 257 988 263
rect 996 257 1052 263
rect 1060 257 1084 263
rect 792 214 840 216
rect 792 206 796 214
rect 806 206 812 214
rect 820 206 826 214
rect 836 206 840 214
rect 792 204 840 206
rect 180 197 220 203
rect 228 197 668 203
rect 676 197 684 203
rect 420 157 956 163
rect 964 157 1004 163
rect 148 137 348 143
rect 660 137 956 143
rect 996 137 1068 143
rect 932 97 956 103
rect 344 14 392 16
rect 344 6 348 14
rect 358 6 364 14
rect 372 6 378 14
rect 388 6 392 14
rect 344 4 392 6
<< m4contact >>
rect 796 1006 798 1014
rect 798 1006 804 1014
rect 812 1006 820 1014
rect 828 1006 834 1014
rect 834 1006 836 1014
rect 348 806 350 814
rect 350 806 356 814
rect 364 806 372 814
rect 380 806 386 814
rect 386 806 388 814
rect 588 716 596 724
rect 940 656 948 664
rect 796 606 798 614
rect 798 606 804 614
rect 812 606 820 614
rect 828 606 834 614
rect 834 606 836 614
rect 588 516 596 524
rect 348 406 350 414
rect 350 406 356 414
rect 364 406 372 414
rect 380 406 386 414
rect 386 406 388 414
rect 940 276 948 284
rect 796 206 798 214
rect 798 206 804 214
rect 812 206 820 214
rect 828 206 834 214
rect 834 206 836 214
rect 348 6 350 14
rect 350 6 356 14
rect 364 6 372 14
rect 380 6 386 14
rect 386 6 388 14
<< metal4 >>
rect 344 814 392 1020
rect 344 806 348 814
rect 356 806 364 814
rect 372 806 380 814
rect 388 806 392 814
rect 344 414 392 806
rect 792 1014 840 1020
rect 792 1006 796 1014
rect 804 1006 812 1014
rect 820 1006 828 1014
rect 836 1006 840 1014
rect 586 724 598 726
rect 586 716 588 724
rect 596 716 598 724
rect 586 524 598 716
rect 586 516 588 524
rect 596 516 598 524
rect 586 514 598 516
rect 792 614 840 1006
rect 792 606 796 614
rect 804 606 812 614
rect 820 606 828 614
rect 836 606 840 614
rect 344 406 348 414
rect 356 406 364 414
rect 372 406 380 414
rect 388 406 392 414
rect 344 14 392 406
rect 344 6 348 14
rect 356 6 364 14
rect 372 6 380 14
rect 388 6 392 14
rect 344 0 392 6
rect 792 214 840 606
rect 938 664 950 666
rect 938 656 940 664
rect 948 656 950 664
rect 938 284 950 656
rect 938 276 940 284
rect 948 276 950 284
rect 938 274 950 276
rect 792 206 796 214
rect 804 206 812 214
rect 820 206 828 214
rect 836 206 840 214
rect 792 0 840 206
use DFFSR  DFFSR_7
timestamp 1733888598
transform 1 0 8 0 -1 210
box -4 -6 356 206
use FILL  FILL_0_0_0
timestamp 1733888598
transform -1 0 376 0 -1 210
box -4 -6 20 206
use INVX4  INVX4_1
timestamp 1733888598
transform 1 0 8 0 1 210
box -4 -6 52 206
use DFFSR  DFFSR_6
timestamp 1733888598
transform 1 0 56 0 1 210
box -4 -6 356 206
use FILL  FILL_0_0_1
timestamp 1733888598
transform -1 0 392 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_2
timestamp 1733888598
transform -1 0 408 0 -1 210
box -4 -6 20 206
use XNOR2X1  XNOR2X1_3
timestamp 1733888598
transform -1 0 520 0 -1 210
box -4 -6 116 206
use DFFSR  DFFSR_8
timestamp 1733888598
transform 1 0 520 0 -1 210
box -4 -6 356 206
use FILL  FILL_1_0_0
timestamp 1733888598
transform -1 0 424 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_1
timestamp 1733888598
transform -1 0 440 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_2
timestamp 1733888598
transform -1 0 456 0 1 210
box -4 -6 20 206
use NOR2X1  NOR2X1_8
timestamp 1733888598
transform -1 0 504 0 1 210
box -4 -6 52 206
use DFFSR  DFFSR_4
timestamp 1733888598
transform 1 0 504 0 1 210
box -4 -6 356 206
use FILL  FILL_1_1_1
timestamp 1733888598
transform -1 0 888 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1_0
timestamp 1733888598
transform -1 0 872 0 1 210
box -4 -6 20 206
use FILL  FILL_0_1_0
timestamp 1733888598
transform 1 0 872 0 -1 210
box -4 -6 20 206
use NAND3X1  NAND3X1_3
timestamp 1733888598
transform -1 0 968 0 1 210
box -4 -6 68 206
use FILL  FILL_1_1_2
timestamp 1733888598
transform -1 0 904 0 1 210
box -4 -6 20 206
use INVX1  INVX1_1
timestamp 1733888598
transform 1 0 920 0 -1 210
box -4 -6 36 206
use FILL  FILL_0_1_2
timestamp 1733888598
transform 1 0 904 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_1
timestamp 1733888598
transform 1 0 888 0 -1 210
box -4 -6 20 206
use BUFX2  BUFX2_7
timestamp 1733888598
transform 1 0 1000 0 1 210
box -4 -6 52 206
use INVX1  INVX1_4
timestamp 1733888598
transform -1 0 1000 0 1 210
box -4 -6 36 206
use INVX1  INVX1_3
timestamp 1733888598
transform 1 0 1000 0 -1 210
box -4 -6 36 206
use NAND2X1  NAND2X1_4
timestamp 1733888598
transform -1 0 1000 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_8
timestamp 1733888598
transform 1 0 1048 0 1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_1
timestamp 1733888598
transform 1 0 1032 0 -1 210
box -4 -6 68 206
use FILL  FILL_1_1
timestamp 1733888598
transform -1 0 1112 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_1
timestamp 1733888598
transform 1 0 1096 0 1 210
box -4 -6 20 206
use DFFSR  DFFSR_5
timestamp 1733888598
transform 1 0 8 0 -1 610
box -4 -6 356 206
use FILL  FILL_2_0_0
timestamp 1733888598
transform -1 0 376 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_1
timestamp 1733888598
transform -1 0 392 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_2
timestamp 1733888598
transform -1 0 408 0 -1 610
box -4 -6 20 206
use XNOR2X1  XNOR2X1_2
timestamp 1733888598
transform -1 0 520 0 -1 610
box -4 -6 116 206
use AOI21X1  AOI21X1_2
timestamp 1733888598
transform -1 0 584 0 -1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_7
timestamp 1733888598
transform -1 0 632 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_3
timestamp 1733888598
transform -1 0 680 0 -1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_6
timestamp 1733888598
transform 1 0 680 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_2
timestamp 1733888598
transform 1 0 728 0 -1 610
box -4 -6 36 206
use FILL  FILL_2_1_2
timestamp 1733888598
transform -1 0 808 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_1
timestamp 1733888598
transform -1 0 792 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_0
timestamp 1733888598
transform -1 0 776 0 -1 610
box -4 -6 20 206
use NAND3X1  NAND3X1_2
timestamp 1733888598
transform -1 0 920 0 -1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_5
timestamp 1733888598
transform -1 0 856 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_6
timestamp 1733888598
transform 1 0 920 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_2
timestamp 1733888598
transform 1 0 1016 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_5
timestamp 1733888598
transform 1 0 968 0 -1 610
box -4 -6 52 206
use FILL  FILL_3_2
timestamp 1733888598
transform -1 0 1096 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_1
timestamp 1733888598
transform -1 0 1080 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_3
timestamp 1733888598
transform -1 0 1112 0 -1 610
box -4 -6 20 206
use DFFSR  DFFSR_1
timestamp 1733888598
transform -1 0 360 0 1 610
box -4 -6 356 206
use FILL  FILL_3_0_0
timestamp 1733888598
transform 1 0 360 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_1
timestamp 1733888598
transform 1 0 376 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_2
timestamp 1733888598
transform 1 0 392 0 1 610
box -4 -6 20 206
use DFFSR  DFFSR_3
timestamp 1733888598
transform 1 0 408 0 1 610
box -4 -6 356 206
use FILL  FILL_3_1_0
timestamp 1733888598
transform 1 0 760 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_1
timestamp 1733888598
transform 1 0 776 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_2
timestamp 1733888598
transform 1 0 792 0 1 610
box -4 -6 20 206
use NOR2X1  NOR2X1_4
timestamp 1733888598
transform 1 0 808 0 1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_3
timestamp 1733888598
transform 1 0 856 0 1 610
box -4 -6 52 206
use NOR3X1  NOR3X1_1
timestamp 1733888598
transform 1 0 904 0 1 610
box -4 -6 132 206
use BUFX2  BUFX2_4
timestamp 1733888598
transform 1 0 1032 0 1 610
box -4 -6 52 206
use FILL  FILL_4_1
timestamp 1733888598
transform 1 0 1080 0 1 610
box -4 -6 20 206
use FILL  FILL_4_2
timestamp 1733888598
transform 1 0 1096 0 1 610
box -4 -6 20 206
use AND2X2  AND2X2_1
timestamp 1733888598
transform 1 0 8 0 -1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_1
timestamp 1733888598
transform -1 0 120 0 -1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_2
timestamp 1733888598
transform 1 0 120 0 -1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_1
timestamp 1733888598
transform 1 0 168 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_1
timestamp 1733888598
transform 1 0 216 0 -1 1010
box -4 -6 52 206
use FILL  FILL_4_0_0
timestamp 1733888598
transform 1 0 264 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_0_1
timestamp 1733888598
transform 1 0 280 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_0_2
timestamp 1733888598
transform 1 0 296 0 -1 1010
box -4 -6 20 206
use DFFSR  DFFSR_2
timestamp 1733888598
transform 1 0 312 0 -1 1010
box -4 -6 356 206
use XNOR2X1  XNOR2X1_1
timestamp 1733888598
transform -1 0 776 0 -1 1010
box -4 -6 116 206
use FILL  FILL_4_1_0
timestamp 1733888598
transform -1 0 792 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_1_1
timestamp 1733888598
transform -1 0 808 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_1_2
timestamp 1733888598
transform -1 0 824 0 -1 1010
box -4 -6 20 206
use AOI21X1  AOI21X1_1
timestamp 1733888598
transform -1 0 888 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_1
timestamp 1733888598
transform 1 0 888 0 -1 1010
box -4 -6 68 206
use AND2X2  AND2X2_2
timestamp 1733888598
transform -1 0 1016 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_2
timestamp 1733888598
transform -1 0 1064 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_3
timestamp 1733888598
transform 1 0 1064 0 -1 1010
box -4 -6 52 206
<< labels >>
flabel metal4 s 344 0 392 24 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal4 s 792 0 840 24 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal3 s -19 897 -13 903 7 FreeSans 24 0 0 0 enable
port 2 nsew
flabel metal3 s -19 317 -13 323 7 FreeSans 24 0 0 0 clk
port 3 nsew
flabel metal3 s -19 277 -13 283 7 FreeSans 24 0 0 0 reset
port 4 nsew
flabel metal3 s 1133 977 1139 983 3 FreeSans 24 90 0 0 out0
port 5 nsew
flabel metal3 s 1133 937 1139 943 3 FreeSans 24 0 0 0 out1
port 6 nsew
flabel metal3 s 1133 897 1139 903 3 FreeSans 24 0 0 0 out2
port 7 nsew
flabel metal3 s 1133 697 1139 703 3 FreeSans 24 0 0 0 out3
port 8 nsew
flabel metal3 s 1133 537 1139 543 3 FreeSans 24 0 0 0 out4
port 9 nsew
flabel metal3 s 1133 497 1139 503 3 FreeSans 24 0 0 0 out5
port 10 nsew
flabel metal3 s 1133 337 1139 343 3 FreeSans 24 0 0 0 out6
port 11 nsew
flabel metal3 s 1133 297 1139 303 3 FreeSans 24 0 0 0 out7
port 12 nsew
<< end >>
